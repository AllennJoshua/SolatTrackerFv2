PK   �]'U[?C8Gi  �0    cirkitFile.json�ے$��%�+#ѯi)����q8K��ݙn�^�y K\�J�LVFmdT�9����n7�hxTwr�Ӭ
�c�
(�P�������i��N�6=|�t����?���{�ҽ�����ϟ���Oz�~���K�\=�����n���oN�8�c?������Ǫ]W������ڌ�I�����C9�f#��fs�"��as�"��es�"���,��.	�?�|�e��xң��07��v��檟M[�a���8t]���w�Y���]5׶��M��.Tڎ�j{m����ȫ�������ڵ�i�j��Q��T]UP}c����irl�S��m�������U��S;T�quիQU.̍5��R���5�:5��"�S`s�"�S���EPɔ�C`\���Q�F6Dd������䦮���+�U]9��Ug�j��镫]8���~z;�<_F.Dd���l�Ȃ�q����!"��eC����!�SX�,�;�3�p���;m6�yR�kO�mO��6|�͆�,�~�Y��6"���m6Dd���lu�|�͆�,��e6Dd���l����������4"���N6Dd���l�Ȃ�;���w�!"��dC��"�w�!"��dCD|�Ɇ�,���Y�}'"���N6Dd���l�Ȃ�;���w�!"��dC����;���w�!"��dCD|�Ɇ�,���Y�}'"���N6Dd���l�Ȃ�;���w�!ԩ��N6Dd���l�Ȃ�;� HȻ�8�-h���o:mz�+����d�*(�UA�C��8�jN�:<�;�@� `��\v'���S
P9��3n�[��3�S08���?ȹ'���ꉟ���C�|����X�
����κ�
ηU=ճ�]oUo�w��߾3� ~�V�����O�VyS�05�M��W]5ͭ��nL���wf5�Oo8��?}6������Os�VUg�Puޚ��i�ڞ��;S)�Χ7L�;s0"��C��o����p<˞� �+�	��}?w����E�~ք�p�-��L�&͛1��-W ��k3!�$ ��s&6�~6�b?��ʂ���Fe����f���B�g�QJ.��M&����~����P=t�>��������O����ʍ��:�f/1�ʂ�vS˨,�u÷��2��ۺ|�Ά��t������45*�O�KS#��ߧ�!�3ݨ�l|����Fe����t�����45*��KS���B�g�QY�}�^���wQY�}�^���wڭ���)5�q�F=���]Suv����׃�����X(o_c?Ɏ�V��{.��1���G�?b�!����,�#�^r���KΣ���{�yT�c/9�ʂ?b�%�QY�G���<*�����Ge�w�{�y�=Q���KΣ���ν�<*���KΣ���ν�<*���KΣ���ν�<*���KΣ���ν�<*���KΣ���ν�<jN�w�%�QY�}';9o?��n'3o�N�u�澮���
��|�MS��~~	a���Î�D\��<;"~[�AD\��|7".�n��a7��ȁ����E��E�M�"r�"��49p���N
�)���+��t�,��r/S�ʂ�/��U�,�s/a�ʂ�3�F�,�^s/a�ʂ�7�F�,��s/a�ʂ�;�F��+����9�� �3M���K���ν<*���K̠���ν�*���K̠���ν�*���K̠���x��D<�.�Ԁp)+����4�]���i�vPv�.Z?V;���Nc٩��jg��A�i,;urX�V;(;�e�N���je���ԩ�jWc����Xv��`�k��A�i,;u
X�V;(;�e�N-V����ƲK����18�X����y��e�'�
Dzt\�LБɂ_qSzVS������O���=�~���O����"�~���O���}.�~��O���:�~�8�O����E�~�X�O���]Q�~�x�O����\�~���O����h�68����`~i�8t���`~i��z_���?8�0���O�����~���O���\�~���O���,�~���O�����~���O�����@����߲
�{���X~�/U�����,?�j���X~�/UG��?���
���'�=ن��d�Ya贰�b�4s��i�Xzpԃ���R/�~��O����c`��Q���KU�����,?�꽁�G=X~�/U���z��4�_*t��ρ�,?����G=X~�/U���z��4�_�M��`�i0�TU��T�X8�p��Á�,?�*Y���X~�/����?��4�_�
�`�i0�T��8����`~�b+V?�?��4�_�5�`�i0�T%�8����`~��/X?p�����Reb�~���O�����`��'��G����`�i0�T��8����`~�7X?p�����R�p�~���*�,�%S;p,��V�v�ι�|��p� UO�q�_�#����A�����~���%;η.�c��"b}���1p��֥r8n��J�q��N��������Q�>B;(;z-E�-��]�[f�l\�}S�N0͕ZU�B�yk���k��$�|&٩�F�p٩�2�p۩ĤV�̏��=�����D��+;u-�zV;(;z�|8�vPv�
������Q�p��V;(;z�|8�vPv�
�ď�.���!����Wp$~,u�%����#u
g�e��hp@��Q�� �:�G5�Z�x���	�_F-�<�~�0�/��bD?p���QK� �8���˨�X��r`�e�R,���*^�1��0�o]*�l�E����+47H~�R97Hk�ڎ���kX~�'� ���x�/��dD?p���Q{� �z7	��k;�A��kX~�'� ���5,��ړx����_F��<�~�x�/��dD?p���Q{� �x�h��ګ�t�ޔ��_ȥ!���ǒ��c����ʗx���2*_R���+KR��`�eT�,����~��2�W�A�C'Ł�r��<�~���o��7�o闝Sj��T�z�뻦��PW���?̓۾��
Dzp���Q�� o;��Ԕ�|�ʗx��1��$�{�1�_F��<�~���/��eD?��_F��<H6<8���˨|Y���`�eT�,����z��2*_�A�G=X~�/� �����re�<�~���/��eD?p���Q�� �8���˨|Y��`�eT�,����?��2*_�AN���,��ʗx����_F��<�~���/��eD?p���Q�� �8���˨|Y��]� �+K�A��X~�/� ���,��ʗx����_F��<�~���X����'O;r5�<H�Ze��:�8n�Z;จX����j�h��=�o%W���ѪAR��V������\�������df�M�鶮���U��Vaԝ�i�z<�T�\˸ѣ��07��v��檟M[�a���8t�i3;�	���E3���/<ǚ�}������n�����v���6c7���زS�u�:Q]b>BvR�M[{ݵ�Wvj��5��z5�ʅ��&��U�-;���m��!d����!�����$~,u(���h&�c�k@�p���E3�K]�ɇCheG/�I�X��O>B;(;z�L��R�}���A�ыf?�����ʎ^4�:�E3�3ap@��Q4� �:2�&䢔x��!�_F��<�~�0�/�hfD?p���Q4� �8����(�Y��r`�e�,���;��֊S�� ��C,��"�kk�n���ۺ�^E0��Ug�j��镫]�/i�r��<Ȫ68tY�g,n���ԅhp�C.=I�
��K;R��`�e��,����XG=�Ҏx��Q�_F��<�~��/��dD?pԃ�Vzr5�B���]U�QW�uuՍj���VZۡ�ھ;��
Dzp���Q�� �8`��˨ZY��0a�e��,�۞��\������~��W	S�Ӧ7��Zŏ��X��*�v��^�'�x����k������{�����7�߷��;����|?�~�~�e��i��W�V_.Id�]q��8o7ܷ��-���v�}�⼽f��弼a�<p^�/o8/o�/�9/����Yo�::���\W���jX~N�]����-?��Y�ɵ���k��|[�S=���V��=�m�<����ǣ���%�05�M�ͫ���V��k7�æ�7Λ����c��[����g�Ƶ�7uջi�\Ъ����[�;M]��sZ��z���-��b�o54��܆�G�m�;�v��α8�W0{��Q��C|��D��{5����P9=��"�nl�l�V9��b?��H?ߎ�H?��HU��F�ƍ��c���+g����<T��0�.6����@���F���o�Js�ctb%tsf��Wk��ϰ�ϰ����O4bFQ{��y�83E��^Şt��� �����ٜxC|ʛ7&
�n�`�i������m���2Xo�lD�byvƛ����f�ge���7�S�q��o��75H�Ov�T(/�Y���|KtRu���I:k�j0�5�/�T�`�7�#i���#i�e4�o<��\�ߊ�I/�6x��1�RlM���}}܍��@
��F��3�)�ٟ�����.���Mz�v� �qV�`��kŤ�Dt�,+�x3-/e��S���c5tS��6�
Cg"�u��M�����5��ؚ��>C3?���QPV����qЍ�}5�My_�m�э�vnb�2o��D��V�	o�e�3�?�e��73�uc��rvdsŜX(q3ׂ���%s�(u}�(���R1�E<�ÜK)v`s������\N����������X_�޻P��l��[t�|F �s|�a:�<F �s�r�͔��x��@~��x�|��Ѷ���4�0�3�Q�j�g�0��Q�bR)���Rr�H�3�@.�qn�5�q���9g�	����v���a&'��a:��R�'R������QHi�����QH�d?j"gp�o���̏��ҩnԔ������qRZ\�q��q��(�t��	��̏�����&(��q������L(�n%�����}5I��ӂ8�����q�:��q��q��(�s�3�̏;�G!��9j'�w0?�BR��� N�5q�G!EN0?�B��`~�9��8
)r��qR���	��=̏�����0N0?�a~��.��q��q��(�t5�̏{�G!��a�`~���8
)]u���5̏���u�0N0?^��8�x�Xpr��4ύ�ִ����&�͈@m�)���~�+j�<��=�	R#{��L=T�b�sf�W�����)��1:,�U:��GC=oe:��r�QW�げ\�*�55�-����]g ���%�C��n���m��v3��`��	i�[�p9�\�R;E_��s�OH��]�,RA��r!�򊨜@H��"*')���	�D�+�r!��K��dQ9��~�{ '�7����@H��D���x6'�G!�򊨜`~��D���l *'�'dQ9��8!����8!��	�D�+�r��qB6�̏����@H��"*'�'dQ9��8!��	��	�@TN0?��ď^IyE��(��WD���($R^�̏����`~��D���l *'�'dQ9��8!��	��	�@TN0?N��r��qB6u���	�@TN0?N��r��qB6�̏����`~��D���l *'�'dQ9��8!��	��	�@TN0?N��n���8!��	��Q�@��"j}@�^�@���WD����x�$2Q򊈌@@��""#%���D�+"2Q򊈌@@��""#)���"q^�a~��WD��܄�"*'��&�Q9��7!��	�	�@TN0N��r��pB6�̋����`~��D�X��8!���	7��M�a~��D��ㄼ"*'�'dQ9��8!��	��	�@TN0?N��r��qB6��Rn���x�T2��E�j��;��@]%�j���m�@]%�j���u�"�Jp�"\�ɉ��Dt��E����Ջ�*�U�pU�ZD�ZDW	�Z��:5"�6"�Jp�"\�)��Dt��E��S+�k+��W-�U-.��EFK���v<X��BA�P�%v���>cW �L�e"/�Z�m�W��V&�a�eئ�Ame"0�Z�m���V&
a�eئ�Zme"1�Z�m�w��V&a�eئ�sme"2�Z����OX��2a���[^�2q�[-�6�e�h+����2lS~���B;bB[b2q���ˌL\&�V˰M�>2���e"l�۔�$��L\&�V˰M�W2���e"l�۔G&��L\&�V˰M�p2���e"l�۔�'��L\&�V˰Mu�d�d�2�Z�m��&��L\&�V˰Mu�d����D��u���H+��(���d��Ca���h+����2lS}Cme�2�Z�m��(��L\&�V˰M�&e����D�j��n���2q�[-�6����V&.a�eئ:�"�:��L���a���h+����2lS]Yme�2�Z�m��+��L\&�V˰Mu~e�:I&t�L&.s2q����D�j���2q�[-�6Տ��V&.a�eئ:�2���e"l��T�[F[��L���a�ꒋh�e�2�Z�m��.��L\&�V˰Mu�e����D�j��޽��2q�[-�6���V&.a�eئ�d���!T�C&.�2q����D�j��>me�2�Z�m��BF[��L���a����v-��fi�z�-_�Z���%,���L\&�6ݗ"b��D%-�V˰M���حL\&�Vg�%ީ����Qa\�k��u��`��@]%�f�^�ދ�׹�Q��f.��u�\��G��ԛ�Et�\���*�k�Z�fR]%�f�^�G�*�5��*��=]3�8�����*�5��j>*PW	�ٵW�
d.n�u���]{��@��F>*PW	�ٵW�3x��+��)u/r��ͯ�Z ��V(쒉�r���"��	�D���^-�Ej+~��ͯ�Z ��V&a�_{� ��L&�6��j,R[�PL�m~��X�j�ۍګ\���W���L�"H�ͯ�JA&(˭fJA&,a�_{� �� ���ͯ�Z ��V&.a�_{� ��Ж�L\�[ʹ ��L\&�6��j,R[��L�m~��X��2q���ګ�Hme�2���W`����e"l�k��"���*[eˏys���"�]�Eļ"l�k���a�_{�*�L\�[͔*�L\&�6��j,R[��L�m~��X��B�2qYn5�X��2q���ګ����j�Td�2���W`��2q�*[�2qYn5S�2q���ګ�Hme�2���W`���엉�ͯ�Z �<� ���ͯ�Z ��V&.a�_{� ��L\&�6��j,R[��L�m~��X��BG�d��j��Hme�2���W`����e"l�k��"����D���^-�Ej+���ͯ�Z ��V&.a�_{� y2Z&.a�_{� ��L\&�6��j,R[��L�m~��X��2q���ګ�Hme�2���W`��
�����r���"����D���^-�Ej+���ͯ�Z ��V&.a�_{� ��L\�[)�(Bn5�Xde��J��ȚU2qYn5S�2q���ګ�H��`�_{�n'3o�N�u�澮���
��|�MS��i���.�|T��ګ��@]��k�Q�Lg��
�5�s�u�\��Gꚹ���
�U�kv�U�����@]%�f�^%*��Б�
�U�kv�U�����@]%�f�^%*�����
�U�kv�U�����@]%�f�^%*�����
�U�kv�U�^"�ɯ�J��˄\"l�k��"�
�d��j��HmeB/���W`��ʄ_"l�k��"��	�D���^-�Ej+���ͯ�Z ��V&a�_{� ��L8&�v��*��LH&�v��*dSA&*˭�Z ��W���V����R� d��ګTd��j�Td�2���W`��
m���e��L`����e"l�k��"����D���^-�Ej+���]��
I@���rk��"����r��RE���D���^-�Ej+���ͯ�Z ��d�2R�������L_O��鍮�V�r���tW����Ы�d�c�h���8H��``Z��X�6�s�s���4�T�(��n�s�f������6.gy�܍��rVw0ahg�s�vQʹk�j�[�@9����e/g�ЏC=st�g�������c��80g���8���a�=������:tS�����ԸήèaVq:�>t�r�5Up��꩞u�z�z{:l(�^��e�������l�*η�7k*7�(�W]5ͭ��n��/ڳ`���P�h6������Ms�VUg�Puޚ��i�����vz6	���H(�_䂭{5����P9=��B������r�����6��OB9�I(��~��8U��c�`�(���?̓{�eo�&��q��b�셄b���4nԾ�og_9�t1���j��Qc���Ǻ�Pu!��BB9�e���C	s���]���"��Ø�L�A
ʱ.�c]((����kcd=W�ԍ��}ס�T��f�~�ܱ!���9"�8���`tq�Ҷ��k����F�ٸ���<̍5�M���6"��I(�mDB9l#�a�P�H�ޏ��T^�8�a��ٴU�߆��9��u�mDB�G	對H(�mDB9l#�q�v���j=�@��-ݍj���VZۡ�������h�C?7~��n����U:��i�| p!�rQCЍ�}5�M����o�6���ƈ��fs̅�r��M]_{[Wޫ�E���y�V�њ^�څ'.{(	��p�&�X��~��3�������{��~��7��!G�}�0��ٍ}l&=��jv���u1hi�1�6)<+�e������_.�F=Y5��iԃ0=��F �����4�C���y���+�F  u^��0��J/�H=�c\$�k��6�ok��F!���q'���0�BRO��N0��a��N��8�|��9qR:� �����QH)#�	7��M�a~���8
)e.�8�����qRʔ�q��q��(���	�����QH�)�������q�z�[�p­���R`~���8
I=eyb8�����q�z�?�p��q��($��`������QH�)g�	��̏���S61�nM�(����QH�D'�w0?�BJ���8�����qR��������QH�V1'��0?�BJ�X�8�v7qۛ0?�a~��n�q��q��(�t��̏�0?�BJ���8��x��$��(ǂ/-Q򊈌@@��""#X��DF  J^��b���zE���`I� ��x�$2Q򊈌@@��""#)���"q^�a~��D��܄l *'��&dQ9��7!��	�	�@TN0N��r��pB6�̋����`~��D�X��8!��	7��M�a~��D���l *'�'dQ9��8!��	��	�@TN0?N��r��qB6�̏����8̏����`~��D�[I�-���8!��	��	�@TN0?N��r��qB6�̏����`~��D���l �"&̏����`~��D���l *'ܚ8nQ��	�@TN0?N��r��qB6�̏����`~��D���l ��̏����`~��D���l *'�'dQ9�v7qۛ0?N��r��qB6�̏����`~��D���l �9̏����`~�D�+"�hp,8�%��z-�HlJ^���Id����(yEDF  J^���WDd����(yEDF  R^�E�6�m��6!�|�<��u��HyE�[�a�`��D�+"ߢ�s�($R^��f'�G!��ȷ�8��8
��WD���	��QH��"�-�0N0?�B"��o݄q��q)��|�#�̏o!��g�Z����F4��� T-�U�p�c����K�!
Hp�"\c�uq�;D	�Z��:-n{G�u��E����w4*PW	�Z��:-nyG�u��E����w4*PW	�Z��:-nwG�u��E����fw4*PW	�Z��:-nuG�u��E�����@&�a�eئ}m��.��K&��2�����D�j�i_MF[��K���a��e����D�j�i�SF[�(L���a��ke����D�j�i�YF[�hL���a���e����D�j�)@F[��L���a��d6d�2�Z�m�ː�V&.a�eئ�m�vĄ��d�2#���L���a��}d����D�j�)oIF[��L���a��d����D�j�)�LF[��L���a���d����D�j�)�OF[��L���a���$&��e"l��T�MF[��L���a����h+����2lS==m����e�2+�Y��L���a���h+����2lS�Fme�2�Z�m�7)��L\&�V˰Mu3e����D�j������2q�[-�6�1����e"l��T�UF[��L���a����h+����2lS}\me�2�Z�m��+���I2��d2q���˜L\&�V˰Mu�e����D�j��~���2q�[-�6����V&.a�eئz�2���e"l��T�\D[/����2lS}ume�2�Z�m�/��L\&�V˰M��e����D�j��n���2q�[-�6�? ��P��22q���˼L\&�V˰M�A�h+����2lӽ2���e"l��t?���2q�[-�6�3"�m-����2l�})2���e"l��t�2q�[�͖x�Nf'�G�qͮ���
�5���u���]{�z/���}+��j>*P���|T��\�k�R��5s��z3���\�k��u���]{�zǞ���k�[�Dt���]{5����ګD27�Q��Jpͮ�JT sa#����ګ��L��[͔:��	�D���^-�Ej+v��]��L`��ʄ^"l�k��"��	�D���^-�Ej+���ͯ�Z ��V&a�_{� ��L(&�6��j,R[�pL�m~��X��2!���ګ�Hme�2���W`�;2q���ګ�Hme�2���W`��
m���e��L`����e"l�k��"����D���^-�Ej+���ͯ�Z ��V&.a�_{� ��L\&�6��j,R[��L�m~��X��2q���ګ���$��L�m~��X��2q���ګ�Hme�2���W`��
�+��e��L`����e"l�k��"����D���^-�Ej+���ͯ�Z ��V&.a�_{� ��L\&�6��j,R[��L�m~��X����L�m~��X��2q���ګ�Hme�2���W`����e"l�k��"�:J&��V3-�Ej+���ͯ�Z ��V&.a�_{� ��L\&�6��j,R[��L�m~��X��2q���ګ�ȓ�2q���ګ�Hme�2���W`����e"l�k��"����D���^-�Ej+���ͯ�Z ��V�̇L\�[ʹ ��L\&�6��j,R[��L�m~��X��2q���ګ�Hme�2���W`���d�2���W`����e"l�k��"����r���df�M�鶮���U��Vaԝ�i�z<e�^�G�qͮ���
�5���u���]{��@f��G�*�5��*Q���|T��\�k��\��G�*�5��*Q�̅�|T��\�k��\��G�*�5��*Q���|T��\�k��\��G�*�5��*Q�̅�|T��\�k�Rg�2Wn5S�^&�a�_{� ��P�%w�V3-�Ej+z��ͯ�Z ��V&�a�_{� ��L&�6��j,R[�0L�m~��X��2����ګ�Hme�1���W`��ʄd"l�k��"��	�D���^-�E�,��e"l�k��"����D���^-�Ej+�%&��V3-�Ej+���ͯ�Z ��V&.a�_{� ��L\&�6��j,R[��L�m~��X��2q���ګ�Hme�2���W`����e$���O?���<�z�i�]i�t�&;VA�
�:�ǡW��*�ǐ���q�65������>0l0��0��,c�i0���y!(����ژ���c0c�cxcyԱ�'5�*NG|Շ.Tκ�
ηU=ճ�]oUo�{6	尝H(��4:���-��r���x�U���|��q8�"���P�h6������Ms�VUg�Puޚ��i�����H(�_DB9�"lݫ�T�����AW}���Φo���#�~	�E���sJ�z��Qϱ�]�C��׃����BB9ԅ�r�	�PӸQ�~���}�L��hj�y�F�ujW�BB9ԅ�r�	�X�q4f�%̽�Vt�������w�S���X
ʱ.��1�vm���j���r���:4��ی��O��P�g������ԃ�r8��]�|e�6z��E�����an�	mh�:n#�a�Pۈ�r�F$��6"���������q��\��i�6�a�q�9t�q�Pۈ�r�F$��6"��	帍T;��U�c �Ɩ�F5WM_+��І�ЏH(�m4���?VC7�q��*���Bu�4F>��P�DЍ�}5�M����o�6����M��̄���r<ǜ������W�L��Y��U���5�r���.��x�KA9�G$�����������p�����i�����p��O���ϟ�aO��������?���K��8X����x����L5��E��
�8W�<�0k=�ϻ�I�������>{lۮ��P���߷�9��U�L���>~��b��׷�P�}����h�v����u1"k�1�6)�=�����zۯ���VF{������̆g�:�շ����(��������v�{�V��[��5����z�{=��i��3L�y�0��PW0U`v���M��zbm�ͮG��`�}��Q7lXo��x�]'��7�u����nG��c�}s�A��d�����8ėo�2������lu��y��n��l�^���Y�o�Y��������5��oΫ���뉁�2�WG�8L�I�P�`¯Jɠ�,��,ɒ���M#��n%C2�����dTf��澟�g����~ƽ?c�6�.m2;�	�!x/��Mb�AK�b~�Iر��/V��^b"fE�t���~��`�v���ƣB�co�b\U���Q�(�d*"Gٷ~y��r��av� ��58���'{L�#j�ᎂL��Ǆ��o��%�� F%��Q���	��5����%,n�`BG]-wR�K%�6].��&�V���X&y}�Kg˵R�a���Zf��֢���={f�A��Z{�NQ������]ñ���._y��5���*4�U��ǩ{��o���g�MbQ�.�šb�T4I��^�B"�a ���m�I+^�6�G�`�rk�}G���G<�ZE��%�34��(���i���d��WN�X�$���8L��mH � �}3�#�d�T�C��=����l��u殺�J�>��}��v�W};���s����x؍�K����hg�B�.4��GC�1,�y��l㛉��HJ�o�I7�ʛ�0�̉��nۿ��gP�@�j3��{�F�X+��i�������`�wY{G�A% �gh�x~�/�H%��~7�r/ɭ ��t@�*���Fr�[2�qc���'ⶼ`o�kLmtBb�!�*חp�0����T���XT�����NՄ%zfoR�p��6�}�n�L��tTX2k�1�����,��ѓ�����)-�8�Y�����]��]'f�R+�24�pr(��tCsC궼���wƙ�m�ԉ�fy���F�o��S��Λ���`�Jv�u��doR�FC��p}S#b�c�w�uTfwѴ,�7	��2ba�����=�\���cd ޴��~��H���j�EN�������[{����V[}�J��*[�
�ݼ�*Ę��}f8�/�/)`2�ވ�	�L���x�����*]~�����%XՀx��ƛ��^�HZ����L֛k��_o���������kC�"^�G��!ަ����:Vp5�F�C���#�V J5�s$�*¢�i��f��=����f��~�ѳ
*�%�_.�y�~���i<u_Ƶk�yƇ����{�7�g�ȫ�跺$�pW�;��Ex���q)�'��b�<������*���;��vJ�[I��үX��ߴ ��p	@�����% 	�-L �˘ , w2X �f� ��`��	�p_���N�$�9�aHr�C�$	�T+�H��-�D`�0
Db�<uĐ�*SMA,��c ��֩�b���5�V@�c ��o��]G��{�
p�"���s)���N�L�Om���ٷ�~@�'��2N 	��� ��9$�7t�I�/��s����� ��`��V|�K<��Eɛ�Qp�'D	�͞|!�|�r��=�|B��>W��[?�/�����!a>�[�Ѿ�kJ!^�[)���R�ݥצ}cw���o��b�[\�z�A����W��,��(��vWv�H����?[�[6z��p���W��	n��%q�r!V�{r������3oӆK?����`\��U�|F�����ܸW!�Gy���a9a���i �d�K����@��%���m��u���Ŕ�W�	W�ie�zÉ�j�q�J��q�Q��Q!��-B����mH(�ɑ)���?�b��Jvfx<�w=��}������gf��Y7�{��.&�۩zhI=rH�= ��0�w�_G����󽚹�ϊa�:5��W�߾/�{������@X�稿�Y� QfE͖�{��fCQSB	[E���j57�;�FeQ\w�l��� ����ݯXB�m�*T|g6���Y��8���R@s=.���pk_w8Ǻ���^��mv�ö&!����r��׺�(�������ܻ���i�}�gĵ����MF��:����;2�=y��v�!������Nz���Y�1or���H�@Vѡ*�"f�nQ�j��v9@��H��^4/ 2 |ۆ��u%��~� ��+�N��H0�L4G'��}x�	�m�M��Ƹ�v�t���7�|Hn�x����dr1��R�r�D)��9�����e�9&�D]UE�zd�x���d2�mQ��	��A����σ�U~�7���u/��wN���g�oq#�Y)&v���J|		;�E,����kw�d����Ȏ��7JX��p�PzC�k�������#Y�:u�5+�]l�i�9��>"��eD ���j�;?��0�)*d�*�^%��U��Q���}�o=�o%]˼�>+��D�ys4!����+#Yz�dl	Ϊ�#ɺ�f�F��X+��Z!�0���Q���η�$�A^��+rT�z�j�KB�vI�K�͖W��Jq�6����e��Q���̃��*
���ȣ�E�V�����Z�+;�C�'�jT��ƚІV�Ñ@�ޏ��T^�9:�0W�lڪs��dǡ�#�Y
X��n��p��L���py�꧷�Y�u,�&�U؄�%�n~p'kk�6gd����/��9�hkv߾>j�:�[؉p1�lG��4��o}�&k����&-��������9�or�����0T�5�~��l����h��=�oop���Xn=)1���uo.I���G8\���m �)ե�/F����"�L>OHv�k0���ִ��~�_Y�?��V-���	ǯ�}K9���U!�j�[���6˿{�n�D�f�F8��e��6���N��f�' ��f]��t�����I����'![�D�A���y��ނ�j�<1sj�gL�{KY�ʭ�Z[���0t֍�o2�#��ESdcf���J�3��8��X��ҢK����FA,����7Õ�T�fˠR�Qfz�n��(v��L��j�C7tU�G]�62�F5WM_+��ІQm&|��df���ۺrs_W�z[�Qw>����s�����ֵ���o#����[��[�'�nߧ��K����xٗ� "M2�@#�N�Ϝ��m�(�!V`��B���G��lv��o�،�c�a�kЍ�}5�M�����8�GS�ܸ��7�:M}��Ə��M��mt���n��n�uMA�=���Cz&���ZD��$NB�x��R�6�Y[������u彊�����]�*;Z�+W���5��:Nb��q����7`mm"���ȘI [��T�YY���=}t��Zio,�Mwb3�w'6#���ng̷�̔���֔(��e�Y���zN���]��/��ܟ�>v�������<?���x���x���8�S��[�dC�i�"H|l��7�f��Hq�w��?fkI���}���w�.8n-7�Wͯ7s�g���Y/I�6ԩ�bC�S�`C�S�g��Pi������X|1#ݝ�p�z�=�3�'H.-���y �,#�Q � �V�|�� x ܫ�W>���t��� &���/�����c�/�G�,�����c���y ��x[>���3������c�/�⇰ ok�Y>F�p�|���� p���5 #R � �S�|���O�����1� �< ���)#� �S>F��|���O�����1"�?�cD �ǈ< ���y �)#� �S>�:y�?�cD �ǈ< ���y �)#� �S>F��|���O�����1"�?�cD ��P��O��.9���� ��A���')���Zn�3�:��K=��$Ž �O�,I1���dDRvI�Y`qoX#��#�3I�qDR���:B���A$���P����DR͒T�#�7I��Mm%I퍋DR����xЏ����ȅ��V�:�	w@�WjqG@�c�+��U�V��Pi�$�&-�s�c��Py�1RL��/< ^��q�bB���8H1��!�j?��c%M�9�驪Pib���*6�����XISaz���*-���M�� x���*���M�� x���*���M�� o��B���8H1�� ����*�{�M��`c��Py ��nz���Py ��nz�����/�;�8����zP�� ޖ�q��B���#T o��<B���#T o��<B���#T o��<B���#T ���<Bݰ ����*�?�M�� ����*�?�M�� ����*�?�M�� ����*�?�M�� ����*�?�M����n�����GP�����E��p�,��)&D����,��I$Dl���"6�~��b?/�Ȃ��Bd����� �`C�zP��{"�'��&sPy <�n�����kPy ��nn�����VPy <�nn�����VPy ��nn�����VP'` ���A偘�"&� ��LA��	T ��=A���T ��=A���T ��=A���-������*�2�4���[\��ă����7� � �a�i0?u�`�,X?,?槮��D�A����`~����y�~X~��e��[�����a�-�pfo֯�����)��`���4��:�`�Z�~X~�O-bf��Wg5��W�	��]�P@���d��X7��]���8�P�����X�P���"���x�P���.����P��]:����P��F�����P���Q�����P�./��b4D1`��w`b���Q��F3L;�h�a��F3L� h��)�t�b�q�A�)`��0ea�5D�)`��0e��5D�)`��py�:�!:N3L�;h�q
��F3LYGh�q
��F3LSh�q
��F3L�v��"�8�P��ZAh�q
��F3T�c4D�)`��;���*��L0x*؂����c��Xtf��S�,���(�P���_h�Q��F3L����0C�f����5DG1`��0U�Ck��b�5�a*k�С�0C�f�j�5DG1`��0�Dk��b�5�a�}����j4�T��!��:Nq�8š�0C�f��e�5D�)`��0��Dk��S�5�a�S����j4�Tc�!:N3�h��>,XC��S�5�a�m����j4�T��!:N3�h���0ZCt�f��S=d���8�P��Z�h�'��G��q�G�)��j4�TC�!:N3�h���7ZCt�f��S�r���(��(�c*�[���
�G�5S�ŀ���`+��[���	ka©V�Ar�@�yd	����ȝ,�/�R`>D?r��ǃ��Q)�zg�~����������Z�����u��|,݌:��;��r���������˨#����/�� �� �~���=D`���2���A���˨#H�^�BA>D?,��:���%�
��A���˨#H���zY>�|���, �hR�Q
�_ FCtdf�S)� �!:3̩X �����T
, �h�K�s* b4D�&`�9� W����"S@G+����^�^mM.���(�*�T������!�aN��@̢7:�3̩2X ����T, �h�}A�8�~��1�aN��@����0��` FCt�f�Se� �!:�3̩2X ��Ԁ�T, �h�ކY2�
St�B/�GU`��J���I<AG1�
��tf�S�� �!:�3̩AX ��ŀ�, �hOCG1�~��Q��Z���A��~K/�GU Ԁ�, \=��t ΩAHU ��+�Q?��� , �h��q�sj b4D�ŀ�� , �d|��0Ü���Q�aN�@���(�0�a FCtf�S�� �!�:��W�+ �h�[�sj b4D�)`�95 1��0Ü���q
�aN�@���8�0�a �d%:N3̩AX ������ , �h��S�sj b4D�)`�95 1��0Ü������q
��_ FCt�f�S�� �!:N3̩AX ������ , �h��S��$���+ �4)��X�����b�J�iV�eN�@<�������S��*�(��u;��xSu��+7�u��Uu��l��O+5�RH�j����f�$�ǃȹ�`Wrn�lˇ��I��x9�*zn��|x�����|<��䵄|<�~X~%	��K^G�ǃ��Q�����5�|<�~X~%	��K^?�ǃ��Q����䵃|<�~X~%	��K^7�ǃ��Q�����5�|<�~X~%	��_��?�$!u�P�sJ b4�G%谄^� �!:3�)IX �����$, �h�I�sJ b4D�%`�9%	 1�C0Ü�����	��Z�A  FCt�f�VV�j�ukK� #):j3̩2X ����vJ����(�^t�� :�����~2:�3�):X ������b�%�
 1��0Ü����Q�aN��@���(�p����̇5��� �*�j�sj b4D5`�95 1��0Ü�����wStPsPtp�����/ӗ�So:mz�+����d�*(�UA�C��8�j>Y��\�`� ��֠�4\��	�vd�אא��p-Q/ܗjpj	pf��b��G�%;À��p��,�8��5�v	Ws�x��<o�/���--YqW��2���Җ�{�o��aVq��>t�r�5Up��꩞u�z�z��W6���Һ�G�[qS�Fg�UqƦ��Tn4Q<��j�[���8k���G�X�cg�Z��4W.hUufU等������>vï���K������`*S�C������*vckgӷ��'3��I�ߙ��~�3_!�~g��9�F=Nը��Q�.��Q]?8_~������Jco8ܲ�-n���ǚƍ��c�}�L�ňn�y�F�ujWghG��kG��kG���n����
s���]���"�nb+u�S&G;
\�v��(pt��ڵ�i�j���r�h��M���6c7����|��+bm�T(p{!��+�p�,�MvkK�[N���4��^w�������Q���&��Uj��H��ςIp;mG�=��Hp+m�1� ���N�ޏ��T^�8��\��i�6�a�qF=t�^ۑ~��o�$���#���v$���ۘ���2�N���]U�1�?m4�nTs��u�vhèV�����eSڍn8���?VC7�1\it��D���n� 1�#��٩!�F��٦��}շs���h�&Σ浱z�	���M]_{[Wޫ����c@0wU��hM�\��
;�����nc�&�-gnc&A�[�Y��n�φ�����i<=ޟ"�׻�vGYi���w��R���=[�M������ٯ��=�q�c;ʹ�\��.�"����"�����������p�ꝇ��<�Fw^Y������DZ=�ΤQ�ŏ(��G�0��GI��CJȳ�C�|������)3���Z�܆��~�2���u�{3F[�b[��֪k��tԤ7��u���C|����6�P�Gקڮ�';U���i�96������Ժ���)O�K��ʸ��6D�UOONCc|�N�Ԛ>�c�?�Y5�x�V��ӓ�v�b5C�1a�:7�f{�G�t?��'��k�[���ߣ8�6u5����ҡ���ۦW��=~n�5!6y�[G�g�V'��E�� ���2�sc���M{Dg���>ZM5�h�n�z�c3T��:���T���0 k�$a���eغ�Ź�[ӏѻ���T�L�ɧ���R]�'�����jL�b��ﻇ�Z�D�-	i!�#�W!�#dVY!�#dW�B��N�8�c;��L�/v�C���rm=GGU���}�7���5-<S��o�e�15�c8�z�a�6��[�p�<76�$�o	��.ҭjY⦋���6Bv��:gy��%�I�X4��L�;�^x��WY�K-wH��%D18n|+W�����2��d�+|.=1�<�z�da�%������Ƞ����k4����K���K��I���*��5���S]NJ\�"��t���,���ϭpڜ5RA���
'��[��:�{�0p�*/��ۍY'q[����I�`������حb�'w����S�>�8n���,-A�� �Ij��K/M�n���ћ4Ѣ�G-�9��%M��t�&Z�ot|b�('���������zCb�*'����6M';�x)J˜�^�a}�5�r�W����kZr����>O�M��$qr�X����R��MbN'���S��g[�e�eu�9ILKr5��&�#f6.�m.ڔ�t��-�m�ӄ8�Y��uc/�[�Te�1s�89p�5�*G+8n�V�iQ<v��Am����X�Kj-�m� �X���vn+'���ؙ#�����C֊���y��������)-D]���1=���ƫ���?������O��Ov�'��'�����_��~�S��S���f�������S���v�'��'/�Y�|�^~�~�h��j�BR/Y��zIӼp1K.�EI��R��M/�f^d6K�͋�f)�y�����f�^�6K���٥�闿������ھ|�]��������˷���o��o0/<͒����,�ż|�Y���v�Ӿ�K����첍�-٥-��v�ӽ�έ������fv��{��-5s/\�����������}�2ߟ>���<+��6�C�߇_�S�}u�}�w�<͏�D�Gg��.b�P�~��y��p���~���q\>�����u�2}���1Dd�_���jR��@A���U/���Sۨ�/?�߆n�ɻ�vq�gi�
��ԢN.�Io��+�.(�>�U�;c9���'oj��r�0T��fu���qԪ�^�pm*�n^�ķ��W�iϑ��DZ]���e�S�������_�+*��e`S��nKM��|��:��������!R:���V��y����=��ۿ���??��<=<~�R�~�qB�������@eL�Q7�F�|��>4m�1:qt�Ls�c��7��]Ո����*h=V6�q�F�^��3>}���}�~C:�����S��=Q����%������yz��?D��{-���w�n��C|��s��W�"^K�3��g�%^��mH��+�����\ �4<�ix���V�%\}��sK�[niU��-�j���U�?�����V�j���U�?����ǖV���Ҫ֟[Z��sK�Z}nŪ֟[Z��Ϯ�z���_�O��:=|}�k��������'����U^���!�+��m����k��!�A�j�4T�kǪ�z���uqx��tǵk&�v��I��c���_�hud�ՋU.������A�����MV�tF��l$迉�������,Q~��ea�A:�F��u_k�Z�j���?�7�d��9���s�Y��C�ct&A�'S�_kC?�t�ɥ��)�5�������Owڏ�Z;�)�k�'���]��.zXh�\��#�f��v񘎳FEA[>�o��thRon������ܵ�1�jL�LZW]l[��j⬠mz?����s���ꩧ�����z���_<�2_+ ��(]g_���+�/z���*�d��J�X�0��E��Wa��Ҩ�����4
2^x��i}��s/���}q|����1�kQ�� �����6]��?O�*3����~T��)���E}���?/}_��_�.�Y��U�������`��A�˨��(!�՛`�]��cє�y6,S/�����)���O@^�Z?G�!Nč��1�.<�P/��:����#Ж雬{iLn#�h7����2͵dֿ4���{�y�����&B��z�[����yn��E�Bxi�g�����]vA���H�㋛�\/4^��,���/{����/{�2p�eT�z�6��Qm���R�Ww���駨b������_>}I	Y_���?�<���ߺϿ�����˗O�ww�=L��/���v��Lg�y��|����տyFNGϿ�~���_��K|��w?�i���E��ϟ~�����?�ק�?���>�(��������/���?�?�"����3߾����?������n��򵗼<��k�.|ڍ����X?Y�>�����|�?�*�����m"�����_b�}�/�c���+ϣ��hB�¶V��ֆs��>���|��8{�x��v}�m���t�b�lU��mj�3*RY���[vD�#~�7툭9/}4N��1�HsM^O$��y_=�~��{��Dg��(���ho�B����k��i�l��Ie��QO��������;�wF�~4�	6�����D���d���#�e�NIe��]O�>A��߶'z��4�Si:��}0�~���M��nZ�r�"����ߧ�����E�1�n�z�B�M�Eۘ��Q*����=.�J��������}��~�o�mk>�qj�:�m�6��8e�>�A*��˧�ʼ�#~��~�o�����6(k�j���]�Mml���u��R������S��������hM��Zg�M;�);'��.����G�����B=񧟿�����o
.������_?}���6�O����/s7<��0=���c�h���_�>Ʈ�r�3[���CsΌj?�8#q��T���4�Ʀ�a�\��6��][�f���k��� ʥ �|Y�]J?tWI�)���c�c�k.����5k5�g����s�M�5ҕ4sqW)��9���t���+�}����J�vH���l�$�I9��s-���:��K���`C�����V���B�8r��܏U;�C"��}3��wu��q$��Eb!�bba8��s�t:�������}p��鳃�`]�tDs�/)��$@Ox�H���>�Ͻ��>��]�^�wG�g��.%�*o����i|�s�)�÷��Pǟ����k|J��$ɿ_����/���?O���4�??L����O�_�W�2_ӑ��1�A�V���?�ip�:�ǻ�]�{���/�8��Ĺ-�7}Wв/�9c=t��Cz��_�*�{2͓{���\��Ö���g�����K���i���9;ȯ���������~s�о΍MO|X}�~�����ǻ�G��l�������X�ؕ5���`����6p�go�l�l�ؠ�5p:lLh��ǈ�5)z7�6��k`�n`S���ԃ�#6�Ranp;`k�v��e\�zp]ԃ��Z�����K}
ڗʒ޾T���^�[�f֛׾�������o��:���;���'�쾽pL���R|C{1����s%���]6���'�������o�&ڕ�r~+c\ʠ�4�M�T����c$�E�Zy�B�n7��B4:�,�BRa)���1����ԵH������[�>0]?�6F��)ẋ��.z��L�&�`c�$gC��W��7�#_�A5{`�6�7F��=���b�|Q+l�wg.��%�`Cf3��E�S�<��`ӮȖkߌ ;�*3��l^[�~r���b.ټdw�A�ټ�~�ra��X*|Fr���6̥O�[����A�3��B����7e��v�K��N�4to�A�ټ��\�&�����$o�|n�\�\�с+p{E�^4z{��`�&���n�O*�x��y�,-�tS�a�Q#4g���,.yJ�<ך3�l*x̬/�_�t���2��73�v��8jO2��c�Ƒ!�m��{���{�%�����N�`���bSlV2�{d,;+˚Ӗ4˼~,\O���T�^�'w�N�t��cٜaڢ�s�[�@'��M�0}ظE�P����\L"����=V7�Ʊ�D,{_�A�of�ޕqC2��c�Ƒ?p��TlhH4�3�"s�n��o��K23j��$���3�Ya��#�j\=��Z�eX�1���[P��M��F��(;pe��LW��9�0��MN<�'�]�>�Wr6�nޠ���c�,:�ٴ9I(t����4��l$�c�w�9/�i���oPj{R�d���X���$�g���V��*w��I{̷�]�6�1��C)�x6F�29���Gi�S]fz-my�-Z�j�ܷ��׼�\�p�6e��eϩ�y����^��|���z�>}�]�9�Tz�����ع�z{��1�7- �?�$�u�WW-��5�-�x�E�o_�e��"V�����E��gZ���Z�:����b_��|D�jU�#H�8����u��`�ϵ���Xy�	7sq�����k�P��x� ��s���+O5�m�fJ�}��=�#F�%w.=�.\��:<WRъ�Y]���ם�TM�&�8ږ\e��c��S��Ie*���hn~\-ԋ\���z=qƖ<������b�L�5aԻ:<��!��>A9��/�W�S����L�Ƨ�C��a&���`��fn\�x�Wm�C� '3���GJ�:�OQD��U4�,2u���z�eY<�c�z |���c��8H�/73�v��86��.�w�'J��#C3�Ȓj�eM@J�3���e��F������rk�#�g�rH>�0!��jD)ڃ]8���y���kc���%4� ��G�wef=\Y���c ���6��Y�J���F���e���vq��r��C�l(٬�V�,ެe����Kl�.�X��j=n�Q�i�^-U��Zy�A��j�[,k[�^"P%���M+H�2��Pŏ
�����9Ry�sfc�fQ��b^��8N�����@������2M��K<��e ���y3�RDM=��BC���s"���I;�Jj�����P�����u�/��W/�?�Q�~�^b��,!�4�kP�܃l ��sCkx�s[�tl� ��X�e��U�<[�`G"����9���Y� �C����
64�x����5�\��Gӈ+��4	]7rI�k�X�X�"V�s-�9��V�� ݺB��D9r���Au �� �����oLڣ�<�xQ����SUוǮ��.��"�ۘF�we�����~�Ƒ����Ϊ`�C�]��r�d��5p�%�I�E��QC�������jL]��漨�D}��r��Ǯ|��1�q���G�we�F����~<o#�H0tߕgYnЮޯ&��K���
u;����eu[Wn��*Xo�0�·ح�z��h�%�*�z��f���_kw6���؆څ�j>�-My��X4���1�Ր�4�jt��dPZ�
[��C0	�C�vsQ'H�nH �nJ�|3�톿�{i7��JHmڍ{�����jf�"��o��c�s��n6��������)6�mt��D���nc�8�/�F��f�˵o��V�Ʒ��8�p���C��n�C��C7tU�G]�6��nTs�����mՍ�"��M͢��~�?�Qx�tJ��[�M{��Lx�<��-�P��V���[3�hʠ��%Ew�h��Up���i}��"���l#� �Ƞv[è�0��z����;�օ`辉O��z���5���M]_{[Wޫ(�i��3sW�ʎ����H��HZ�EW�]��͵��>����8����l{iW��T�Z�*肇���5�%�x�-�QW�����$��$��WV�ZŪi���$�[H�F���4�JZ=�b�͞]��[�>��)����ē8T���E?�à���Fin_���5�q�"e��ī�I-Rr�&��zW�U����{��2���_/�{5q�=���'����]������{�8=|�>��!����?|�?��߻/�t����O��8��5}������PK   @'U��8nx;  �~  /   images/21dc82dc-72ec-4a9d-931e-ac94256341be.jpg�gTS]��C�"
HMQ��[*]�J�ބ ��"EzQ"]���"H�^"] �HH�u�3�x><�1��័̵3����X{��wF�'a	�����
�@ ��� ,�R�s� mm�6   @�[7�֠+ �:  �o���m3�ە�N ��> E�;@~�Ns^6 zU����Ѕ.t�]�B��������ɥ��q��:y�<�DE�D�DEDDE�D��e$��^b"bbr"�r"�\"2r""r� @�L�����=��߶Hj��6��4 ������'��O�By���^d.�Ѕ.t�����9ې��<7D��m�"�3� ;aH���W ��oA7��s����u������_���������w�O�,p� ##'#� ''�����a�����a�r�����������'���s�������;"�`~YE1!q	��*QRR�P�0��2�q�s��o��	�S ��� �Ӄ� �������������SPRQ�;�]>����������<XP��� 	=�nQe���V�<���R�)x�Vw1�@�[{�SR1]cfa�~�����R�2�r���kh>|dhd������������������@ċȨ蘗��i�^�g���zWPX���CI駚ں��Ʀ��޾��σ_F��'&�~N�,� ���oln���cNN���8���2.��HH�I���D���=	)�(�e}r��Wy��(��WwQ���=~P1�I,_G��ߑ���?��߁�'����|��P`||���۹�A���7�~�^��d[��NŮ�D2j8��;�oD΄�c��-�}V��+�6.��%�:���t�X2;�K�M���%l�q7�+:�i#��ῠ!yp�7�pT��� �H�# k�l�r*V� �D�C�"����O1��Z�ydI��lv�Sҋ  �t��ϴu 6Gi�=�{��7�:V�&d	@q1`UA'���]�}���Tl!��)^E��W���:��h�;�e��&dvq��/K��'���P9o�qL4�[@����y[[z���.oE+����!"h���[��( ���{�9ļ\���m�˅S�z0uhE `��?���xٱa5GI��0�x{�G`��D����N ��p¶�1��]%�����3��ʐtW/�rO@QB��b03��!�R	��% *�Qu�^�'��K��0I
ۧ��a�2��A|�Q
_�E ��B3�S�ՙ�N|{��,[�j��ty��*�e�*n<Yz���AQ��$ B���l�%;�������Z|6�.����;��N,���h>�Lz���	q��Zt��e��9�W���a^͇wk6�ԻË���Qe+P�9���Uw�_t�&��to�/dY�t��פ��W������#-�&3N�M)����J�A�����f�4���Ţ[Ǒ {@�ŵd^�X �-'�v��s	;�#f>P(�6�4�D�ܠl�����,0�%J^'Q2�9��E�SQrD[d~�#��I��>"�K�v�K�e2]A�Z��
e�/��kB�Rs��3b�e:&��%$�T�������� ��~���7QQ�H��?��x5?�v�a�}A�P�F��H����D (^�Oq��� ����%'̿�DM�T�h��:�1س��]�s_c,k.p��ӷXb�QS����wC8:P��}�'�-�l��գ�c��F/�SM��V����Am��ީH�/r<-��*��i�)��@���zRw����؝ ����?��x�*���Y����XG*_�� �g�'3�n�Q�_�W�/��t�9%�rk�$��L�_X& �,���kP!�Gv��?�~�ShW����h��JS�#����]4>�!v4\�f�8�{�suW��a��"|Z�3�(��4���j�1Te84���|TI����AgQ�Һ�6��[�@PB����]�p�.�n]�x5�y�,c1;{�u�nVs<|�tR)������M�^���1��M�:�����O	�W��Tx~�>Y��z��t��݂�EV6��n/���LG��o�D�#��:x�����K�a4@A�'�@c��h���T���(�ϏYt�Q���?,�-V-���tl���=.L��֒�Y�h �k
�*�({#�����Ms�f��cmg|J�5"'Y4c~�qFL�����|Ie����LM_��7R����I�e�>aea�V�%� b�0 /���q��(�R�f%�8����rOi�v�0ۅ����8�1�5]�����"T'�'�O�J*){n}j�Ye��"�g�6���rJA�ve��B$M�3pWP�.��I��X�h]`�-2��`5mP�%R^*�iS�TUܿS���-�+�g�7�-�z��p}��`�`K��J�Kv��AM|�o@�F����8�,6"^~��(Eh$$�aq��U�Ity����19����vz��#�A8sZ�2�g�R���6y:�t�ϏJ�W[����u��F��̪iʒ�c�	��kH{�Nt9�������[��+k�r]�s9��g�č��e!��t�DR�>���y���d�����'Ka�~��L��2�Mܷ9Y\Ynߛv��t�⎄��>�)9o��~M�|o J��"�O����~J�/�<�u���i�>�����a��.���V��D�M���N�S�M��*j0q��o��Y��u���އ�ߡ�{��O��l�q䁍���g�1.���9�V`)2����6��%���E��E����hS��0���9�?�M�U!�%�w���v��L�Kt\O�\�ʪD�Z�MO���O:'�̏Ns�:��燊6l��r���xb��a�b��6'���Lޚ��-?�e���'���D��m$�����-'&{�2K�'A��<��-z2�����H	X�����CG:O��βa[F��D�1��2�,�U��o�g�wnG�E>���=��'�]����"�������X���!f���;��3I��F���S�Z��\��������6�K��7���&�.U��ښbՉ�4��j}��Td�1�i��2פ3�Y:Ċ���k��n>�d��WT��͓��-�Ȋ�P�W�_hp��U�?�@��X�P<nݑx8O�[�1X�i��'��t����Z���l�@�(LY
!�e-S@�4U6�Nf��},��m�l�ޯ�\�W�EVx;��_}����E�����bSc��z�.7i�QJ�f�RGv.������g�H61�=P�����q=r%����N������a�>Kʣ�ۙT��� �g@���l�y�S�ݢxi��Q��3ʔA*3����#d�%+{��Y��ul�u?˵��`�y�m?�S0~@"�Q4h���^��j�Rw2�q܁*'7�����@I���m����+�)�g��/�t�9<�|�ޖ}0r�_���w�~lAm�d��ڠ��Y��41��q�A�Ҫ�����+�~��+��ٞԏ����.}�Pu: �ԥ���~�}��[��;�q����W{��;�}(��d�=zL���کNv�O�Tɂ�^qnZ�`��sS�u��LF��xFvЉ�`�WEQ�>.���ZP�M�X�`ȳ�2[N(�,� �kF�e]X����0�N�E`ߵ;�@��[���cv�8��M������O�>G��,J��T��|a�J|6Yq��^�f�4�e�� ��1"߉<�Ds��5S�"{��z����I����\*�>K��<==Zi�64�6�SB�P�Q�3�}��W]�T069�C��_�s��ȗ}7l��p�?���x���.*�6�1�)r{x�S�c�>�盩�{:�-��>�/2{�Lr�EC5L�B�Q�I2ǜ�c���9S�޴w�uX�f�&)ik���`���c��L�s4	������Wt��2�e�Kz66�}��gS<�~���d�Z|�Z@��v/�R���5vw���c�O�wS0�JT�$o���"��DgS��Ԍ�Ԍ�8�ޔ�r[̞�NM��9��k3�Ӷ	��5�[T1�?u���ݧ��]6BWd?���#$GL�,�%�f,v��v2G
	Kp�`JƀXQ����?�{J��3i�}����,ğ�fu�?j����a�OE�H�j����~!W�N��d͙��*\6�}/��&3;.���o�z$�4�U�<U�H<>��/ٿw�!�{�ؑs��)w��g�P	�����(S��oR�3�s39����{��~�����|^6�7��t!?�1�z7�N��{L|�w��~$;��f��R�,�Hvo��P���[y�)3��pߙq�S�����e���Ew��
0a+����7�M�Z馰��bF��"Aμ �&�^�Ё����w���Z�5�J�;V�zSz���Fy���n��w�ǎ�]s�9�#A����yz��aC�zDz��0%�5�<�-Q]C>��:���Uʫ,������y�z��<�w��'�_�*.�l��%��T��1����L����yg��\k�{�9�>��ct��"�z�-�U�4u�� qTTq�V����N�O���ػQ�:ሢ`j�s.n^�R�\RM����2���`�y��v��K����gH��8<m�)l�����zjo�-��Z=ו��ꚼ�Q��޼��"h��e�=Ԙ��"d��]�M���W���+�j!{������)�2z2.��8�V����k��F�e/W�Q�1o)�k����Ռ�{Z�����봎��p��C��\���)��^ o� P%��*�ߚN�B	��S�'�������^��x����������[x��~ISB>����� ޝs�}�����H�]�`���ʥB���Y&Nn-��)�=�z=SMOf��a�/$u�뫹�n�/Q�A�ʝ�ש-�ӄe�G//w9aa7O!+[�����U���]XTHDP���[ٸ�yqY�98�)��t�s9�*�Kj�h�߳stR�{���&��F֖
��R��suw����s}��)���w�r��_��y 
��r�U��q^R��g[|}}�|Ņ`¢����"b�bb�����n^V~�n����ྜྷ������̍믲�5��K�����V���^���VR��J�VPT��J��V\T�V\�VZRTF�^Ԛ�_tu�7���s޹��=;+/��#���������걻������������������v�������?������?�~��t��\@. ���r��\@. ���r��\@. ���r��\@. ���r��\@. ���r��\@. ����N��Ն���"�/?��z&�DD=�Er�$��keR*rr2
*j*jj�KW.�^��DM}��2�UFFF�k�L�W�^τ�|RJRRJZjZ��m�c=�'��� ���L�����p�N�W�nE-�Y�YC�H��t^촠�ؒ���gN�|��+ %�DЮ�I�1�Mtd�<(��#I����c���nxq�/8p%rrƔ����W��+�eyY9����Q>��̑ع��#��S��!j�"�թ�(�����q=��v��1q�����Rۼ��{x���BC^��|0�h�e��bˍv��p�i�YAAT�g�5��<b�Bqis��@�zL-A h7v��$>]o�R��P8�k��n�� �8֪5��։����z�e���o��Ldⶎ2�w���D�	Ǚ��hni���g���Ζ(�o�Ř�����/�
֥!S�n��:�uN���Z����˪��E���7{=Iw�g�����`A0��9��=t�o�Os����'�p�& ]�8�>>i�n�]~P������fS�؍7`}aC4��6R�9pw�v�5��Ġ��V�+��Y�}�}6�C���PHf��:��ބ��8�^�i<�0�����"�`G��VK4or(9�s"ղe�6�����d�j�X'�U�i�6�J��,Nx�ot����S]D�C�����ow��j�[��EcO����6țh<-zw���� ���b���+�3�b(�S�G�p:���eN�j��� ��`�>�uX��GhN�9T��_#�}
���!z�sb�8B��B�&Y:�n���d����Ǌ}r������ë�o�h������uTU�p�7�tۛ�UG�z1N�������%eA���$@�; �����r��f�^Qnx��Q˳�\��ȁ|��ĿoN2�[�Ο�*J\�|�?E :�y�Ϋ2��9�*������Y���l��rB�m���?p�Ձp���w��_W	�g���{���O �Yφ���>�y�k�|���KJJ5���<�>���j�
7��4ۡZl0�����No����tle%,4�\�;�8A�xE�ӎ����N>p�}��r��(0�/�~% �SCv���5�X�S<'7V� ���'������
��l0i�snw��y8���,�|�j��l(^R�|H��j}`�k���&MX�CU��[�t��Ϡ�!�9G߼�{'�ҫ�!�Gc�pמ�ѥu�ht��c�����6q�a�,�&����M �$�sߕ[�x*F�ҥ����'�4�7�1����O�?�vJ>Dr�G>zޥԮ�p:c|�d��m8^Z�@�\<c����!%�#̪�A��{�l����B�q98���k���s{}ӧ�ڡ�a���^��E�'Y��80cC�	@��'+�3[���;{��>S���ʸ�����eN3{ч9`�ڴ���W�����u�	�e7E_��p��hk��6�����6ƚo���H����F��V�ԏm��\f��5��
+�7:l��q8���'ZȾ��#CLB�4���.^����X�#�Y��p��,+�s�psG42���i�l3t�K!`��+t��sF�گ��`C��9x	ܗ�oLW:?�
i�%���#�v�4�~$�#���fz�"gv~��R�JU���KȎ4D�AN��K:=t���!!�Q�����N|�r�$,�!��_��Yhc�p�SG���2��u.'�?s�R��y#�`���+�d�R�	���	ha^/��ӯ���B�fq+�zP\�����Ҧ�Y1R�����1����Duн��~h��rK0����nu���Gy�	��1�� DD+&b�����c3�� ]��!��(n�����E^ѳ?��MV���?���{ԋ[�3Li�x����Q-�L�D[�-��M���S��޳��PD]�q��ULF��B鯑�/c�z��S�$v�V�Ca�G�H��JCCo��3�Jsۧ	�yݖYO'O�/�B��"�	Ԡ��'C}f�]a ����-8��N�L�������j.�1V�o��ˀ�zE���e�
��N��v�g�
�C�X|Χ�V�Vƃ���L�R8V.޺�S��Lig����i�}2���D��>��(�/?(|l��<��`��gx���P�u6���.�9��PN��zN>x�� T����u_c]�l<���b�*��7�Q�y�̛Â�����c9\�Pe^`�Q�E�`UO���f�f�ߍ����R��R$��{>��z�1Y��_gtsU�|+��g�����(�΍�M|z�C�?�]b�[���	��뙣n�%d(�gї�l,iw�m�Y������r7���Q��n��ρ�|oA'��B���)yA:�Y�2��I���n0�󢲏nM�6+͇�7L7a�2�ϧ�a�j�#S�6�<��r�#����K�ի���X.�T^~���'� ԫO�,
t^|�_}l�d�2��F�Am�a��ϦN9�^z������Bө��Y�?(�&#�̩H9���I��rm���>T1�MS�V��
�%K_�KW��དྷ
�9x6F�Ҵ9$�0��й�>z)�q}2��� )�0��K�]9��`�V�*�+��9�����}NV?O@t���C�ο��\�[tJ��Ѝy�#o�m����8A�θ �#�S�Y=s�8l鸽=�=}��[������d�-�	��va-4F~���ca"V�4�NfIB%�O7y���8���杶�n�t��d�
&��"��cVdp�zKc��(�f����j�mݖOJ���-�m�~��q�Z��|^�rWъ�Eq.���c��m`�}x��մ6�cK�V��[�V�ef~��?�������c�O�������k�c;R��kѺBq�\OM�	����͑��+�vR6|��@3y�ذ�$�C�7j�?k0&Tq��\��D�.�u��hӳH	��[>ST������ڞ��V;�8*�8�u���<���E���r�^�J���j���YZ2HM׋O74L�վ��8w��s�-�+�<ℕ���]�쬗a���rɯ��X��&8E�5�����vd��<�(��7꼲k}��|���&~��G!0I��Q|�&,��	���v���e�Y8�j�R��١@�+ ��m����4�jB���yY�iPU�r
&jU��3�}|�Us�5�\U��窑���U�eW����d�_���Z;-���'a]��8���X#Obgy3��7�ED��D�MេG1h��/7��{�����W;�����9]iZs��, 'xׄ���q427 ��ɕ�D�+\�瞊=���f�?�qͺ���z}����L2�xol���A�?��7��Ɓ`�b�Ԏ�oa��/&���Q6Azucv�.�c��A'#� �6��l���箰+[(��f�^�<�]e]�x�w�,��Y(�Aݨ�iY��ᯚ��}�*Y��Z��:��<& ?��Z���nd���S�/��S�y2�ܘ��S�����e#�t�}j��G���*ә�k-a|�zۢ�/̿�<h>��;�=hY�Z�zqh��#�'\�'� ���7m�2�H����)q°!�~�'�!/[;�w.k��*_7���K29�b�NM�as��;Q4����J�/�.*�)n�8^{��(!H��Pq-F��C}��c��/Iv��!GE%H�EI&�w�<Y��'ʬ�_��4���[�.�V��s'��)?ޮH��7�ɶ���%&��sp�����A�sAGkc4�\���9��R��ڐ�|u��4��v���)*5����j���
��%+QP-��Ϫ]Ssϡcͱ�r��P)�>YK�d�����12U�ϧ�:�1���2S���,�t�%�#@*�*�sC%�]vt�,���Ą.�]�~�O�q��}ݘU��pr���v�ʌ�x_��G�XʧDQ�x��W�^��R��:�{{-�e���EP�B�c��m0��87��z�y���s��'��;�]��
8��?*i���҆,*�J�%^�lQd��h���|����/Լ7��?P�˗�ǌVo�e�l�w�� ������H-5I־$����R� �[2�aU�!��"���������2a:�孬1%n���$6.��B�&r���\����c���Z�OB�u�-U���2q(����f�x+��G����{����S�f7w������ʪ��:�CD����0�+��Vx��V���v�u��?�u�E�A��Jq�~�l���E�ݾ%`?d�ކ�ñ�8�z��'̺~�&꨺Q�_��D�W�"�@d~ߵ��ɿNŞy��z�K/C{nVLiT0i��LO7
®�B�k��:�e������Y����y�]_q0��q���Y�HѾ������	pۆ�(��&hu�r�S��c��t���3�z$�$n��@&Ṉ�8Je+�~fӾϦ�E�[j�-Qi��Z�(�]�6[�*z��[z̟�Ա��A�?�5���6�0C����SIwb��>��f��!�8H�xE4���Bs�Sq��6�����SY��$�	p�J��+L��;�`�j�4�8�H��������2��RI�)1�Mx��~��^usq��(id}�\���G@Hh�u{g3n�h��������g�ں0���ک��L
����iai�7Z�T~�Z������m�;�Z���w~���=���-�u�nn�{�>U���yy�n��	�(8�����F�)�Kׇ/@i�8j������"ä��"�+�ȇ���u~�.�fN<��Ux({����z%A�VU��ѭS�[�j3!��KRg.��gU�N�2������ћ�Yڸ��K��
����w�תRnڂy�X3j���Ǌ(�+N$	]�Cq�Rn��T�%���w�i�$f<b����;B^g�zym�wWM},ž?��bk����?&��ga����_Ɉf���r5���X��C&��P|�W\(n��W�næ�H�eZ����[�v1X����m�?�yƣ
���v��0h۳�O�؍��h&z�^��$/�J�,�����C�(�GN����+�GmӍK	��׳elp7>u������pɳ ��6X�F�HC��D8�q�UF�Q������$��[��k�g���� �J�o0�A[aWo���ZW~���1΅�
�/]���u�x澮��<l���q��h~������'��͘�S"'���ӗ@��b�;�Y ��A'���+H-��a���1g���W��_�a놱�4����JY������d�)�Q�Dq�Yv��YiJ}+V"H�s��@��ǩ!no�W���ry1�g%N��ך�3���G�S~�FM�$K?_c�gW8�<��<��pb ��UX?X_%��D=����e��p���-��|���K��>]�i�F���X1̶渂�O.G]]�y����]#j�5�'ӯҝl�w��.�=�:��CH���U���n��ʴШe��D~��$ۉȻ��O�LN��P:��y�sO�S��:����wi��b(e��(no
OS��� ���х2]p�z��H?����h,�n`^KX���ٝ v��1S�8�F����n®���������b̎sĈ珼́Soqg
�(���P�f������a�^z�z�k�־L��u�/����wĎ�6l��n�w^^��!�������)�q��->"wr�^>T}��Ѝ�A)�s��N���P��D�Y�H ��0XL�n��]���ܵ��^_���2��wvܬ(���~�P2���*~MD>�)4����}�g�$�ҹa�-��j��rg.s��l���?�7�3�k5>�����.�q��k����7tT?���&�P��#�h��=�h�
�DM�T9��.q�J�2�(0���K���~޲���EʦQU
_���$�s��(�F��Z�Z�.�v�4���r�
�5~�}ەh~���L6�1��h8�զ�4�X��h�g:A#���i����@��%�'B)[U��#�YvF�a�_�j;�=�'�;�|)�/_���C��� ��Q � )Ld�
Zd
R)t�b�nv��?�$�08����`��Q�����1�����;�=�-��N��-���q{���4�Xj����͵�͙}Ӓ�5Q��u�5ڃ_S�F��m�[P� E�~��G�.��j�M̼�_�,��4d��}����Gk��-�6���F4�6�'a��!�6G�_�z;�����K� ��ڈ��A�c����zWlf�<(�� �Y�幺ڕ~���k��H����^����;)���4�u�0���=	�?g;�����0K��%�O
�nuZ�`�D|$O��L��A8|�3�/�
H�"�|���.4��n&��-���!�AJ�u0zL��$����Ձ/g����M���?[�!G�3L$Z�w=�:�nE��a;����~�Ʋ��g�g��$�t���O�r���s9�o�sR)��������Z�Y7�INIb�W�"�|ѽ�_�y3SK����`Q�;�������t���d؇f=�[��$��d�%²fo'n��=8����3%�D �_F�spB��O%��2W`Kj`B�ֳϳ�߾�98�\������l�����ol@��(~2
�۠7�A�ba�����l�����ݧ�'�I����$P��R�~�����Ѳ�)Gw^�ӕj��Fḅ���X�7fueqG��q��`��#V�7����d�Ԅ�&N؍�����:b���Y��̱%�����[ٺ'�NO	��PW诇�Y���+jJ�_��*P��Nu�����5
�Osx�Hƪ���w����=��j��(��{�:�����G��k�S����՗8-���F��/���w���hX�=�-O��Ʃ���f��aK�����k	��MBۇ ���tS%5W�@��7�6�Dx2�}2�a���2B���Χ7�2���*L�A�"=C�/��џĎ{D\5�YoS�|	������3��6�y��"�9���T-�)j��xӄ����������	���0�۩���8�oF&�%n�������>�?	�W=7�v55���j����mꚾ�v'�{0���T8(�1ݩ�GE�N��8J'���8K�#�M`��P
dO���9`�q#���䊮���LܶkrS`�/��	sW"��A�v�����/O���eI A�����.��L�i�����i�����q4<"Z�CE��W�+�aV�oc?��R$G�d��_�n}��,�yc_�%@�C>�nL�3.߀ҹ��*17��v�h:���y=.<����{�Ր_��5� W��m�E�+E�V��X|6(T ��a�u&38ӆmk�)1<v�M���ƙ��Ʃƭ$��ߪ6�.�S)2�5��^O�
L�^IK��7-N�1��D#�9��:j�f��v��c��E��?OpG�%R���6_)/�h�:R���ͮ���K�Ѥt��K(]������Jk��T��N�ޑCs���H=�.��w�+5g�8z��6L���v�[�R���S�`�������u�̀��4ts�ۓ��G��f	J��A�k�0|� �U�O��n[׈�Dǅ�I)������y]<KـV�Zj�p����Ȇ��YE�f,f{�R�Jή�c��5tK�wH�˿�hh).C��/S��0E, zs�Y�M��̻[�Y��&v�2�����W�������|]z�T-X�Å	�`R��?Ur���1�^|��K�^���4Ϛf	hk鏭َ�t�a�#����n��:[3��P��8���f]:Mrk|j��2b �޷Js\��M���E'6�oݖU:�Y�F�C$�Jw�h�Z���I`�]!��}��(�x��]�\���2�>��q�(�:�1j8.�m�7�+���79Ο�����d46�n��i6I��W�}#p�\! �z��6��v��U����Eٸ�� k����m$��D�ʎ*~�UC�m��{����"2OU�
痭Q���*劢rr�Iv����S&Q2
�Y{��ޝ|�=)���b=݅f�ъ��_��R5O��g<��j�|\g���|z�:1�;)Ĺr(=���^�w[Ϋ'��؋KT�$�b�H������9AY�0����D�Q�PJr��-w'���\;@2져_iO���D�y��B�x[M�f��/���n��e0BLqv�ҷ���+БDV��735m����(�W�(����bE2�3B�+Tܼ4�jd�m4���q���kaRlb���A��BN]��;+���&�q%)_���FI����%Ȥ]P+֎7 6X��sB)5�����O;ȷ$��,�ុ"��׿Wّ��W���wo��i��z�N�85GGW�Ͼ��{��*T�JO��&�m�3�	}Ǚ��s�~�y�f�↨Ⱦ�����bbE)B��pՖ��\�P�w�P��&���/��hv��I;��������懡����|�yNj���t��]={ʖ�G�u�#4[����y��hy�ɏ��0���e��~�G�.6p<J���s�7I:�RH}>-l��B��������(��!��<���v�}۴�
5	x��Mռ��ա�h�����ʌ�s�I�A^�2��'V�?��ߞ�_�떫��ʹ��A��%˰��.}��ˣU[���ᶜ����/;���mcCE��L?��	�R����T��*v��Vձ�����O� Ap���g�>�)�xch�����q��=S9��\��ؗ[�8K6ʬ����Gq�B�v��.l��f��!�]p���9n�ҷӤ.(N��{��X�e����Z��-���_i6|��j�ڕ���,k����Wc�Oy�+�v�8m���'Q:$ �}y+��S9��m�uC lf�!<r-��0�~ѓ�����-)t2�U��]�)�~��ܤ���f���VN		�.R#y��*�ϓ�k���U � ���b]qT�_U?�h'[�����?c��v1x������]��\�9�G���@�ma�[o�t�T�b2	�-v��Y��"V�>� �`���g��M��1��G�߭S�Հ��d��F�U;���N�������[>�C�u8��w�"�W�?N��۹J ���������'���)���t�ӄ��3~�]u�a[`����ק\��ZO3�[���v;']|���ǭ3�|��!�i��76Z�K�!�-�|N�>���f�LrB������/9G����ժ�GA�q�������G��#��4T~2/��v�W���!�4Sl��z��=0I�WG!�}O3���=��Əm��vs:���8��,U����Ё���%fn�NfI�G�nk/��� �L߇���ɾcx?x�cx����Q��^՚�&t�����t��0����A I>S:^�i����蝓p�8��\�ܖ���eؚ�E5�#W���Mb��c����g!ְ�S! pҐ�S�����в�5��%����a�o� ���m٢9����Y|`���5��! �}!��j-�����k,����[�?	����q�J2�NHAl"V4�N�Smk�u���}��[�S����@ *��"?���+P/���<���Q�3&���+b�)7�8Yk��V���P(a� PK   �K'Uu��@� �� /   images/626defbd-9ffc-44de-b7fd-54699b7076eb.png @迉PNG

   IHDR  �   �   _��/   sRGB ���   gAMA  ���a   	pHYs  �  ��o�d  ��IDATx^���e�u��sz��T��Cu�ht���� &�E�2%�Mky䱖2і�-������Z�d�$D (�ADj4�ι�r�{��9�;��>�VU7��kf�9U�;�������_��Ѡ۳^�g����Ţ1�D#��Qo�h8�����q�B!�'	[8�N�m�5F���FlH6$�E�Q�'̵~��bo��ă��o�F�c�O����Y������>�3ΐ�
�<��3z�7�>s����<�~���^��W$�3�Kq�-
�B���\;&q�>*��x�{�#����塐/�� �~���`�u��v��#��o�+���7
�x9�;TG��s{��\'C�]����3��?���t:�k���L&��G�g�%ߨ�*���yL�8'�u�ep�O�=�и�W�����&�^� ;�[�$x-���r�.��'4��I��^*��M���Gʣ��W�Wݩ�'G��8���uG��z������㱄˰����:�]Nﾧ���c�]�h2��w��ʇ|�������������=�K��������W>'_*� �u�W����q-��L�j^�OE���G���v/_�ޠk�T҆(�X:k�t�c�Pb�[wh�1�Z(!�m8���W
 8���Fͅyb$`�t�]�����1�&ėq�u�������]��y�d��'��jY�V!����yW�F�޶l*e{�����U\*�x��Ea�hE=�!�%��е�];�<�h�����Я�~�����C�Pz��%�)�v�:���5uh'�����P�.��~/�S��t:*��x҉�w<����PV�Y�kS3e�yY�w�A(L}�B��o�ʂӟ#�[��ҡ��gܖ�iC�����В���H�ĉRV���#?A988�#*c��v4�i�#+Ԛ-�Q'h�u�4�h����}�sh�^w�8D������� ��Ƨ���I���t�F�哖Τ,��8]u���^�������Dߥ0�#��u6�廨ן���V���E/��ƭX*�o�ѱj�
��c*��Ig�o�%~P����7�OF_+Nɩ���)�_G"��J']+ϓC�����U�KFpA�Ĝ���8s���ȫ��f��F������_��v�E=d�T�)ψ���@��Q?�Wfff���j�r��'��p0�uy��V��a��o�'�o�{@YC��:m"�)J!R�<՗����_PFte�x���o����@�T]���s�U�o���'�Kr69��䈐?�GyoKG�Hfu�^Uw:�g�)dG:��<(��3A^9��)�sIʣz��C��w��Pz�8�d�����qں���P^�c����s �5#�3J�ȅ�9y_e�F���g�!���D���� ���"�c*������DOx9�����N'#^'!�+�W�y��DE��A�e!*�����=֗��C�!Ⱈ��4`�����_��MƃL_=�J'��L�ƫ����#�Mw�`T��x��~H���%�o��kL5��M�D�r�!E.�G��{1���c$�BŘI�0n�w(M+=�,������{y`N��9�w�?�\EU|�����Q�'������?Ӂ����T�N[�:L�A�A^���L�Y@�A黲�3��N)$�zȀ{:����Yy�?��KA�Q)�#����{�29�-�!�'���~��zc��P�z�EAx��G) ś�g�ذ���Ċ���(r���ؘ���O�#f��wxQ
x\ve��[�	�yә��h���x$�	*@�Q�:��tpy� ��1��F�BD�S�3�L�3�)3�z��x�ʸőѪۑ2���I����i�C��7h!�%��@P��!ũr��u�HD�V3 �:ďz� ��e�\���F�W�U4�̠P��1�R�����(����t����oS
Q��$�k㉢�x��\��Y�V�;me�������"��I�8��O�]4U���y��:I׈/�
��dTW�w��[U�W��*o��dQב�<aq�?����L
���E���3�����m��uH^&[�뀒W����@^T�T 72Q�'Zė��"��]�>u��pTX��N�
	�_�A��k����|'^�܍�8�
 ���?�8�_��Ȅ�:1���Ǌ�	�)Ǹ��������"~%,�� �:vw���<ny>7����N$i�l�:89�6�5I"�٨�/���V�ҥC�k�H���j�ߡ�RE4ЭJ+��
D)svbP�.ޅ2&4dn2*G��d�����ͫ�$֡���buJ"(���PC���Me�B�Ae�pD�!�P.O��܌_omm9*�������
�������QB�#�%��$�� ��ʏ~˃��"��[UD�d���
�T��Dt�o	���h���@U��.
�	%
I��-����ҁ��^�*_��c����K��Ɣ?W��QԷ�n���(�P`�X��'�(���(�զSG�, ��Tn�!~�o\�<����|����t�؜\"�ꦂg��Q��.3 � (_�	! �!���v g��[��"�����Q,��,!
^�j�*�/����5J�������e�F�u\�\͗�7�; 9Ȓw�
�<)R�Z�k�M&#/&�N�z�_���\�Pt���'<�7f��|�h�H��O���9�!P7�Ϋ�kɣn�Z��C��4�8��s>煘d��0�f� }�Wmp�~�	|A=�Y�W�6�e|%����^X�b�fE+�ɻ��<�.x�m��W�\O~�|{�zw�{~�W���yW��A4���C�*���Yy�3՗ʍHy{zʃ
JP=�Z<���lfA6yN:��1�:��ʚ���*(:>�zT���	���]-�[}?�z?�G}��I^ES�U�T����Wv��{C��p��.�w��Cq�U��?qE�N��r�;�P*E�M�����]���	�Uзе�9���2�7�$=uʪ�c�;��+	/�Ho8ꌺ`���_8k���>f�1�%Z�F���P�:m>j@M��r$� !���&�
���R(᰸AMA���\o)d}1a����O��G�Z�wj������tT�1:8�	I�#��!ݾ��]F����nK�Kv�m�pݰo|��đpWZ�\�(jqR�~7@�:�&g/��0r��G`�T
'ď8D�*�뉑Q��'G2F�!�D��1���|�����*R�j����N�"�^���h���=��~??C����#�G R��m��(�@����o�l|D����=)f�e���S	�az���A�Hap26'J��$��;��� ��F� �s���E���� ���1�2H^����7jB��W� ����+hB]�W��ķ�r��$�d���#R5Kv��xS�I���,�J����}���mj��y��|)���sI�9)f�
�b�����\ǜW'�.��n�����&�"��x�����\(�(e�����A�XT@HZGr%�[� y�@�P�d\WMd�yPnG��d^:Ee�{ �c���F�E5�p�kz���J����Q�5~�o�*=#�@�!�������W���y?���Ûb��
�y���Tq�f��6�O1v��{cc~��}���+�w4��.U���׋hť�'�c�յ{�K��t�K����uY,����������E�͝�3���{zW��˲]=��%0��C�x&�»����L<T�6�N��+�D����H��2�F�ĸ�m��_4���ɺn�H$xK!� �z}����	�X.�m!�����C�Q�{i�~��٥V޺����q�����-�9�fe���;ט"�U�@٪BU��\����bPA5A�QЪխǡ�����I�R��j�r���s9���<<fĉPߝ�
!h]�=�
���lo�}
t]�陲����c�����	���J�V1N\e)y��.�^=���+����^��Z^�h��$�b)�y���n���jI|�Ǐ1���(��	C��Qqo���]�ƑgR�T"���w�))�p̸2
�3X�+�j���`���2r�w}9<�Й�3F^&��hA ��@ጀ�*/)��'�d�ȼ�g�F�E;,����W��O^S�����8Swb,o�!ny�R�P�QQ��V�i
x]G���H�*����P�b�kO|/��ʟCq��o���n��x�������i/�@J�k��c⒢��}�̓�-��4$ޚ�OC?�ݾz�[s������(U�gg����Í����uo҄��
�[�[��}`�aϯ�+0�!(�ć\���6."����w����@�����J�.���:�E*�������5�Dd�זb�C�
?�~(���3�Tu�כ��%�
����û\(���@����<�(�|Ҵ=?W�ZǮS8Zͦ�tH�Fu�=�7_��.c��6�-\�\B����@P^��x�B���� T�z���!���dX?ä�C�EiI���V�����Xt(&�T����#c��=9Q�c)NPR����V�U��-�)+��]�N�����d-45G-�p}��o��o��{ߵ����rGl{��ޒ�Od���G)� �	O���C$< 1��^��w5�(�B�z��k�,`LW*��zp%�?�ֵ���PB�SŢ.�2y�����%}��$R)���A�D�L.�!G�"�7���W�O�
��Y,bz�Q� b,��bUl �]&¨�j*s�C�#�[��=��?�Y
Sq�Ŕ_Ϥ��e)b�D����������AH)0�R�2	��CT��Q���S^�ޮ���Nx��Җ��AC�W�+z���<4pB\JCE�rp�κ���ɸuP�	hЗ�6�H�aG9*��ʧݨ��q�l���ȉ+U�j&�XT})��D1(n���ᒷ/C't�{�-�N�w�=+�A�c�X�Ƣa"�Đ��/���:�#����)� X�~�dC�#����Ah���)~�:˻�3!|��ޑ
h�r!�����-��2�@$�yW���sW�z~���#F2��ro�
����3�>
P6�ա< �T�:!�G��?Ԫ5ޅF�+P���{1�].�F^� �~�����~��$�Y|(vO���
���.!�sɤ����&?	7�R����_R0� ����V�RFK�]y��}�ջ�?��X�*>i�����E��u +O$�y�����a�/����8J&|����mz�
,`CyT��G��6���݉���S�r�P|��k����@eQ<��Ґ�G>���8A4s��p/�{=ҙ�x]1~���?�2��"V�5]��\�h���&y�h�UG*�����=�E�� ���Np��$窿p�E��{:ճ_��;���n�i��n��������1�p~ݪ�5�T���2��QLQ"�v��;bDYv)I�-)[@2�n;� � �:K�8���c��]a8����)�b�4�srD��xG�+��{ތCB�ʓ��ꝟ�UC���Q'����8��dA����ȰtoZ�����z��t�����Œ��{8W�md`!��h0��S_��P!#�
|A�t��◾��()�w������	��a5G�"a�V�傕ɤ�͵�R��6���iB�jr(bb���+�����߾�+e$��I���d���m�)��L����ꐼF�qkf4"+E�����TJ�S��0Aܒ�,��Ш�\�;���w� 
�Vr1�Ow��Û�0Zě�脡o�VG�h������yG��K �W���U'p����UoAK��?�QdKu�E�嗧�fG�"��b㥫�5�b�n�.(Se��� �1�䡑>T��a�Td���t������%ߩt������U�|@)�t:�l:���xO��'P�����n$��ԁ�&Р��7񚚵�Gʛb�!P�{�=y��X"�g�B!��M���U�{ndS�4�@N��wm�ZTr��5j5�9)r�g�`��^:��]����U?&ͫ��N��<ݕqS?��$�H�zx�j��t�(ɾ�Q�a���8��U6]O� r��䓻0����3�5��o7�7��sp�8��Cɺ��xWzZO����:O�u����Mҷa1���ĥ��v]���H�ު��g�foxYewPN݈/\�_� Q��	�upE�%��b����U�u�a����p�~�g�݂�����^B{��{��ֱ��e���Z*JB=1J9a�"�*�tFa\I��2��@B�^�B�HF�wZ �"�Nl1�8R�Ba�Ԥ ����q�� f��F�="a�>Bh��9�ħf;1�Kт���J�H��K�!��Q��ʁ�Q��FR��R5�
5�[�"��2yWy��π�4��G������z7��E	�*J�S�!��sU��o4�1J!�ve$p��B�z_��ɋʯ�JWt��2xQ�֓���裸�N�tT�u���� Rr�
��xd��4A��O��Q&���x
�"4���C���|Q&��$�2'FG�Cq)~��x�ʤ2^qbl�m�(����[�@��.o= ؄o��}��7�	� 5�
��x��y5���F�yiZ:IaG-hT�O`����I�0�/(�Lt�&r&��&?�)���v�'��(����P�hN�(/��.�����<W	�2'�(	O��J9j���)Nr�|��(��I�Z�C�J�OK٨Ԛ���AiR�σs�(�y��z�+~���K�%�|��ٗ�Y!X6 �8�XHE1F1���!�𠚐բ@4����(����.���P��$��
 p_<��1 �,�)�jM/��(�>_h���|�r����-���l
�˸.����{j�Qֈ��
�2��Veh�AqG1da�h�ԟ' - �F�+�)���?հ�h���e��S\�Df~�{�\���x5����(�)-�7r���8���ك�b���{ԽF�)�r�Ĥ���s��"�Sy�Qt�Oe�Pz7,�T.^r(L �<�g���YcI�y�-����h��2���?���� �D�$
���(�����2��O��$�:�\А�Cdm�w4P��m��z�)����"GNz(γ�Ǧ��4y~�������7{a;�մ�^9c�aԦ����e�}
���P���W&1��$qdB�GMMR�2VR��\֍��_O�	h$W�,��[Պ�aŞU`{�:Ej�S��!>��C肎a�;�������y���Q0T�ʒ2Ā��O�^ǀ7 C=ҭZ6�wTvmo�3q�]�q�w9��!/#��r�ɿ��56h�0)�:k�ǡ�:
�˳�諉�|�d�)ۀ�@�m<�V�W
�&(ڀ��^�a]}��C�K!���\LBE��ԉ�B�ᠣ�=��&���� �0n��Qq����B��k<�a�C�
F�Y��нY�z}�:(7h�!O*KD&.ӆ��(K�2�P�Q#[մ�e�ŷ��&���A�]��Š`�dХ�%�04�G�n/4�l�ܶVm�fJQ�e�����WQ�"������U��Y2Z��K9�9갲�C�ȣ�|�]|�?K9��C�@-��(�>e���-;����l�V�PB�-kֶ( �*��^d�!���XP���h�&츑�&=j��9��������!�Q�E*N^j�U�Q�=�hV8�^+�'d����s�����:u)�o���d�'M�?S�l�����u�Q�|��Gf�xB��$Pԅo��Q ��������ԣ�0FV̢�j��9c��%zۖ�Y����6?�Ql��ŷ^�dV���f�I
��%�x5�O�M�)�}�|��IS��U��N9����@s�E��1����
E��j�ٓ����l����C�1��'�n���U���}�&D������o~Q_���S~�f0�z���o�8���JV��y���{jQ@�/M-\}�gy*�e�����;�LC�9ާ��+d�8 �B���>�E��=�(ؑ����;�G�Դ*�O�J�L� AN� �চC�#�#������"��8��H(�f3�:a�N��q�T<]�]��)�}��Sg���OT��d:Kw����@�6���S;���'�*��cţ>VԊ�E�u����DĦgK����o��k�8�{˲��=�k�>���R�v����g�J��9�����h�<���m�ܔ�#bV�)Cn�\f�;@!����7�ɣ*��+�)i$Q�TtE/����
�����R�f�b�x��g��)�������+p}7]*��c���2�*Y��G��X(�R.�2iZ��<7gM��à�`���f�@��.���MD���`L4��)�тhS�,��DBG� I�(��(����N��VYF0d���#e#�=S.���f��4�n��0;M�CV��r��a�FiIa�M�0�0e�`Ȁe0���yRT���3�#�:�R)y��Y��Eh[M�@��^��^A+O�A��Tu)ayX�*dH1b�r1o�<��#Tw�2��y�!*�1�:�eL��"�V�S������K��=�#	'y8ݧ2�O��v.���������n��y��/�����Ǭ�~�Ӱ�a�{�~���@��m\:K�e@�&#hC���#֐<d᳚ի��c�H�������f��G�W16@ߦ��#������e	�i�O�A�$H���M�mf�huxeD��o�F�:�q��槦���q�:�B�P��}�V.�0(E���/��M���8e�P�S9<)��.���,}�@:�7�� �� ��~(P�p7�/��Jr��<	�&�@u�W�8^\:�oG����n������h�߸`������f�V�����.ߒyu�(a�)�W�_����JCV�)�2(=񐀖�8��Ϸx(�s޺ �$�S�7�s%5ģTʲF}`@�)���O<���95ʱ��d\-#�U��(�\��:.�
��@�I~�ȿ�B�u��(�ZU��k.�U���d�,iz�O�F�jpGV�"�wTd�Sj�Ѩ���SE�p �#�Yڨ�BeN�[�]�Kn�O��K�s��t���T+�z�>����NZr0.*K�����gs�-��rs�=u	=�4�Tu!#�V���JC�+)��P�[2C|�{�w��~&dR4P���*��:���V���~�b��,\����<ʨ�nn�'����0�c�x�B:�=+"������Sz�.�(��b�a�_ퟚl��-��x|Ӹ�
К�qū�ɢЗ1X��l:39��x���!�Utxgh�ʃ��拶��`3�� U>o*�Ki���9uG�|j�eH}CL�T�q�8����%�>���{UD�wfg�6=��!�?s�al��s���ʲ�&f�ZX��in���d��?K���ͣl�%�2�U9���!���V�<�&���!0��36�1�SP9��eK�O�9h�����ㆃ�5�7jV:Jcff��.#XF��
��dn�l��#���ye�(!�Z�daf�(�R�g� ����U��,�KS�i+ϔ�<[@��5��R�(�dZg���4t �݇)Cco&Fa��[Y�.P�Bφ��D�g�R�%WL��ʬ�3�7`z�!W���C���S�%<E�zд[���/|���3vס)�G!^���A��M�)����SwM���7m�Ũ--�sEM7A�D�g\h�O�����S�4��ޝu���|��Z¶��]����~;�H u��&��L�}+gG�	�g� G�B�r<��SFhS(fm	:�p���ƠS��Є�H����8!#��R��������b���BZ�1dSI�S>�ln&kW�i-� R�İj)k���,G��ʼW�+�0��t��-�lE�8XY�v���\�B��)��Y��O?r�����)��?�}��y{?`�3�����ݲZ�����Ͼ�2�]�����ȑ�O�x��D�|�rbl��Q�Ő�(z"P,�0jݪ�:U��Y:�YdL@M3�C��40���L)m�W��2��[�^}�&=AN��٩�M!�h�F�F>����O�f�K!��C�Gm�����Mdm��͖3 ��� #1<�j����ΣK�g�,�FǠ?d4cKs��S�<�~�Q��2�n�Ik�X�n����m�o�8%x��a�(g�[q�B�h�8g04ew�R���ѳiRn�T�瀾�b�*H���et�ta�z建��!t"2��
9H�i	������ P� p=7��� -v
�Q��<�d��(������"
c`�e�O�\� �3��Y�� ��Я8_ ������x'���>��$0)OT���P*誶k��R
�G⸐��	��h��\]��(*�CDZa�MA����5�sn���R��~F� E1�ެ�����-I��Z��V[ۮ�@ �p�jtg�����W��U�V���d�p�K?B�-X?���Wk�Ɂ���j�J���5��o��E�u�&�Q�è5I���%�B0]�
��L��[�;��G�!�hAס\��.�j'��j7����T�?(3p�+��5�O�7��8Q� 	1�AE��-"٩��3T;7��0bm�J��B�Q8���Vmi��&pk��`ɰ~[ͨf�[� 憸�XZ��[�vi @�� �:�s�	;�y�P�.B�P$IY��jk'�6��h4�Dо�.L5�5(����ۈ�������B�G�{#��J�jM�u��d0n(�(�0�"0 y�[߁wՠ�R����l�j��7[���� ���X>�����>i��p�|�%@�,�$�ۆuu�g�U9g��7-��ӧ��P�����;�ʞmn4\a����iP{<	���`���p�7����g>f�G����K��m
�O�C5db�_���h�Bȏ�j6���+��Ja`�� . $��L��ऄ1�H>ڹd���f�Mi�._9g�L�V1���e޵(ƿ0��tn�x��=�qiڢ�]kU��*E0P��HXq`uE1|�x�}��o|�Dq��[V�cY��đ_T���l�ͤBv�Ѭ����?��B����U���\��$q7w,�ٵHk�z��lu6脯[;6��[*�h����oX�}][,^;{vp6k7�u �Y�+��W ���6�aז������m�IcT�[D)�{�@�c�g1h#�J�qf�Tώ-gm �����l�O 	aW��A�\�VG	����Յ�W�HJcJf �jV�"s��!�+����{u�PG-,�Ɋ3t�<J����T�w1ZK� �ᑇGj��#?2d�(��#n8��2��5MjI��Ճ�b`P�|���y=qK��0���k��7/�4�V@2����Z� m!y���������h�<�=��-.��P_������S�`Q���������NB��U�sE/�������N;|d��V�4�}_R;�13��a.�@�zh�<c��������{ �8!Q��x��¹����UM�j�ka@b���jZ�'�ћ45�1�����[��,���.���H�F���4�B󏴖�O%@4�T�����玖�ҠW�Do�������1�TTC#���F}�e�6�.�&��"㨡�"J�޴j��̺��Uy�W�lRQ|���U��K^F���Q�>o�	���"�;<ҲNoUmP.ݫ`�ۭ.�F_��mo%�y*zOt�!��=�>`(�x$!���v��,4�9JE$yʯr`�(�{{���2p?�BO��ղTI�BAk�1�� ��W�B�^�޲��=���9�!���@�5��A�P�d��4$]K�@���ƨP7q H_�D#�BO�"�^�Z�#��@���P��ɜz'������]s�d�Bԭ�K�����C$��S�\ٸB~Z�N�4P@���PSq���;|n�����"�a��O���ً�Шk7[�n;h p�8��q��*��mc$;��*�UBlX
�Q��mgo�u�Ǆ]��k��^����v���+վ��c��[k6Hd,��C�M�x����}�����3(���۱���P|�G��B��m{�4F����T�Ok	��C�4���ow �1�F��>��.
�������l���"���ٴ�9<{�Ùן�N����͕RV.��F���&<Y�.w�m����(x=�,X�Ұ��
�E�8 c��o4P���Y{��@�R+]{�s���jo���t҅$ul�E!����x�[p�v�1�����o�6�u�t�-�O7.�ޱ~�r��lY}�
�^��V{v��7�R�.xI�9�����x�M<e��ŷm�շ׭K�G�6^Pi*�!��͵���߰�3/B��5*��)x��G� $�
�(�ox0�l�t/�j�q����s���Ր�]���ˢc��).``r���E5�O��E�Qi�V���o���P&t�+M��G��<ߺ��-Y�j� 6�D�^�o�/��G��h�����,�Q@���4�	aD�0����6C���܌������:�B�4���-OM;��؂weP+��Z0Ѐ���ˁ=PS(��0X�V#���+Q/AW�t9E��7 ��K�Q��m�ʕ�����Hq,�X̡Ӻ����:D��j"�4�zs/haLm}m�<t=�X�~Mu5��4���7��hжl���G��g1xXE��^˾��Y�kE-_��rj0�C�R�	5�@䤠>;�
���Ġ5�L�%
��2:ʸF�iЊwd�OD��R�h�����=*D��[����s�S�U)����|n�L�vwv�����44]`�"�ω!%���hͶd�DEk,)t9]�7K�լ���x�@�ss�I�#֨9/�!Fo�����3QY��5J	�ۇ�Z�Z�SV4��<��F̭�v�k��jB?1��h�T�>����~
0q����$nU���Rs	 ���]�O4�LC�շ�2�$�I*oS^����+��xIh2�G�s��O�4>�ou��#�R�>�� 
(i
���O�P��7���[��n�&�UF�e S�Շ�P�[*��OL۝0���덞}�[/�������e~*e��X�٢�ߞ������/� ������?�I��n�{���I��n�C�Sv��9;{����s�LѶ7wm��G<	���ŗ����w,�[B>�ޟ�k��� ؿ�7�D,J�\��C�V �݁]��s�����_�;n��_�����������>���`9�ȕ�g1�C�W^y�b�D����������~���g�������>��	o�^�����u�r���O|�����'�S=ix����Cv��E������+��`3�)�O���k#�=����F�Z�]JpD}�}���y;8���u��_�����y��s���Nۥ��øα�}�O۷���uU�xu7����������~�}��c����i�]8����Ň����W�A��s�%;�2e���[�Gf�ˎ���s6�WwG���m�����n��|�N��=+v�Ñ���<�hw�<b'o:d;�hu/o�6/�fI�ϧ?~�=|�vˉ9{���v�-����]:w�6/�vϻ�\�[�O��9�Gz���ߴ�b�n!o�ܸb'n>b5�l@%�=Ƞ?FV�i@<��Ԩ�:����h}K	7):���ظ�DFj �����ѯjl��lj>����.Ɯ��:"����/*A<Z�E�Q�dOFFPT��5H:BK:�ЌFyI��'5?��گ ���-�Q��� �T���!9�V�	x{�/� ���+P�s0��e����+��y�� ~@����\
��[-��y���Ǥ74�E�4�FND��$v� ����#�0�[(fkk���oi��oY��%Zq��"$��v����^;j��e����NA).)wyf��FChM��a{H�e��E{���Q��J�E�QA��R��$����YZOn ���q��a�>_�t�Y�U»qv��շ��e�ǩ<��m�'qC�IF��+��Q��8���Su��W2�o�U����"�Is�dSd5l]si&q����^25yBK���P�#�����F9��񾾋�O_�C��ےG�����B�Piʅ�S����!6��*���a�|�a��������|�6eW�i�Y
E�p�AfQ#�D�JQ���Q$�ʓ/.@���@�>�Y�Vq|�~"&ntU^����4���/G�]�C��w�1�)�&�?����R�x��z���֣�vh1�2o�7��}�W+��O|������C9���p`!g�s9;�Z�R�ڭؕ�
���|����<�?��{�����Oxs�F[N�B���n=���4|�G�ѓ|4���7رK�5�&��*;g�g?y����Nر��-"��-�ɨo�ȁy�ݴӧ^ǩ��`o�_���>y��{;�t�`Gmy!��I+fb�K�nb����m�����#��?��^H��W��Bڎ�����ܴ]�p�.� R��SU��C����Ż	�H<�������-<��o[���)<�]{����ߴA8�����n�^~�"��{��7��J��{�}7�_��?f�w���'m��s;z�hw�|܆����3x�{v7F����C���L�n9>g��<H�����ۭ7���K���gwڢT�����_x���hG�~���ێ�����#v۝��C>�ܓ��u�n8X�_����/����=�p���E�[�GV�ר�峯�q��2������~��n����-���N����}v�G�{�����}n���ॠ+�=5� ���i(�	+�Q7�dC̯g�>B�PPSM4*T2�?7�snC�"P+W����m����~�!�$CFHs�$c�s��	_�H��f׼�ML-I��#�RQ�!ܛ��4:�������zX��W��� ����=A�@�U�j�!/j�(V�eS4�]�G�O-B>����hڙ���2���2�4�����SeG�W�����Y�|O�4�ڃ��`�ţ����82xg�����gl����U\��Pn�V���!� �u_�L��aAo
�!�!�X�Ļ�H�Q4�*���XM��ln$�"1R2]	�TCn�xuhx�b�ћ�V�P(8a5�I#��ޮ9Pb:)kyxZ�Q߄	�PMW�dB�+}�%�d��/�T�o����Uoy���&ջr'��Fy���5�	}h��l�F�i���ʫ|k�)l�Qg���K�h�t�|+��am��K1kt�#��M�g䟆�j��&ժY6��y�S���2\j�j��c�����"���w�">�q�kԱLV�0h��/,��$~�
�`bs�hRi5����� ]�	��U�ĵ��h�yw�KR�����B7��1lY!3��8i�z�?�g�;k1R��4�Y�v4~d�=m[�{��?�E��-�_�K?e�P�q�Nqս��Ԕ��`V�J���h�/\��+�-���>v;�E�7�޾=��e��3�r~`<R�c��V�Ͳ���^�y��+�寿d_}�Uk�q	�`}���-[)���{o��[�jq��L��vpE���v�ԫV·0v�GZB�}d#�?���� �7��^��}����|���'���Ө�\�s
�c������o���c n#����sX�:��.yT�����9����T&m'���Go��n��>��G쑏���矅}kT6�c�e?����B�f�KR�j�Ѵ�����c�>����`���\��;!t��"���/Ȗ<����=�J٪v��9��#�د`�O'-��MQѨI�XC]_ޫ��O?c�D�>��[�g>q����4E&�)u*�}��<�[���oۍG���6��؉���C>�G�׮T��ۓϞ��MuOL�(�7 +@Կ-�&]�#7��.�����R��Z�4oR+��r^�qҖ�k�"���S z�+l�L#�40��2ԡ�FW��)�zK��.��aS��������4t�� �&�^����'�&�3�)�B��(yP+T�R	��y Rw�� "�j��mH#��c��>&��K�v0�ҋ��I�|�.D�KB�e��ۨF��h�C���4�*P��x�=L�׮e�MO�p�0x�xx���M�4#������w�@�����m�ʜ]<�[�{�hYyzFk�q�ѲN�Bp��5+{0ODذ�ϐ�<���]�n��JJ�7�4S����xh��3>ܿ���ʿQ���t�IY�VG3ą��!���0;k<�.���M�r����jB��Tə��gJE�C�u!㹼4O~zV��GF�"�0ͩ��6120R�)߱�gͭm�X�����5bL���bw��_G�5��n��3����q��oY����R�\*�Fᷫ�4	m��a�4WL�ki�>�bP50b�[�QF�`[�iT�VnQ�c�0P��#���Ug.��_hX{�Q�:��<9�5m��/-�IX����kZ���W�&��
&a5��١�F\���ckF��7�����0��:eӰ��׮U|�_��\ȫ�T�*��������Ԛ6W�E;h^ �����Y��mR��ٶ��Y6_�����q�n�q����=lsEx��=����+����ūN#���ˏ�w�|��:�g�/Tlq�="�����Ϝ���|oo���v��4l���A~��W��M���qP(�_>e[k��;�X��j�7�o��l_��s�÷��5i�~�2���.�jC���+/��_�c{�oZ!���8i��8e��v��yr��k�t�F���}�7��������zԖ�5��mI��vm�~������p��e��?�����K6ҝ�Q;��釳��'���7�N�:F��k*L�TS�&j��5����`�:�Kv��VΦ���м�uˢ���ì7A.#�d/Ү��K?n޲l3�Uݸl�����SoW�J��K�zv������sv��;~�G>67��7?�e{��M����KifA;��vO�;�����O|��a	�е+g޶���}��'�[�|̾��bO���%JK����a{��g>���O=d�$�``ͽ��z�
�3�����x��݈�׮Tl��uˍ�@,�!�2��������?��~�v����D�%��	�d��MtF*�5�c
���Mmj�UN�Q��@��0�Z�#�E�Q�Fy�з5Ů�g40P]Ce�������i)���y��S��iK=Kj8+�~nld5�V�m��gp|�,z` �~ �~T���Sk��_5C:e��NΏ�M��?m�#'��Ä^}�]+�(��h���/�Ad�E��k2��0�_�5'��Ԋ&�[`NY'�ZyG�
��U�=�feL5_od�se�$3�����ѕ�ܹjG��phD��tUG�ch� �Y��.,,�`���=h���� HY�)O��&���	�������Z�!NJ6F�91>F$���<���ׁ���5��W?�9��r9�2���\kyR����'����c���cĝ��
1�]C��(��2Ϥ��P��0�W'�<Z�9��5s���xٴM��#'OM�9)e����9Si 夘Z�"K D�<h9,����FM�q��ޞ�dkx�Fd͔A��3��(#^NL+�C��ʐ��9M�Ф�*�o��CAuk>������xYj�����m��X����:嗇�!.�_nݪ����v�o��	�=��v�����C���>�ɻ��O�i�~�v���{?y��|����lv���*QhC��Dh��TQsk��(��rσ�@�4�P '�ЫI-�r����)�8�l�4�)h�Hy��(��XH�fv,�ߵ��>fs L�&�� [�a#���u��ן����o�o�_��b��~���ڙ��ux�B�$���C/����._Z�>�7�V�b4/��vê�i�Ө9ya~~+،F�!#����'Q��}��d�?n��>{�}�;N�A]��@^n���{�<��s5%��O��i{�{o�o�Ο����7H�E��{N��'�[�z��^�-����mw�u'4,��c���yNZV��f
9��ϣ�hj-f����tuț8t�7}��p��� $--�h�H�b���b�����ٿ����+��y�tc�b�`K36���D(���,!���<�V&7�$�������ݯ������}�����+g<?��e`���CKs�/C�K���o����������g�g�ߐ��G��=��,�{u���my*a�hSq��������?�����������T�A��M�;8-�%&QA>�������|�N�ڷ�]^���<d[`;?�G_`���^� E����6*b�S�M`P�t ����f�[�z�Z����y�)H�˲S��t!��M�+���`�M�Z04�7a�� .���U4�d�^u'D;�DН�>�����ޕ�Vپ����a~���Ј�"�0�t���%|�6��\W}���� �L�SӼ�Nm��M�Kw��4�y�\��}M����S�O��Zk�r �z5S-_��ֶL6�W����ao����Kn��(�L~��W*�R&ѫ�n���Th�� N�B�Z�i����D�4j���Q��IMj��zvj��Y�,!WT�B'e<-=W���)P;J��YUJEF��R�Wj�<����*jw!!��×�0���z�ʃvb� "/o��֮㹹FWM��L@%(5��}�2JRD��}��iI�iT�-���X.w�HF0i�j �rޖW潉�7!U%b��e�@$0r	�/A�3��sj�H>EK�L�y}��Sh�d�
Ω鴁כ��<u��KbPeʡ�{�
�0���5wfP�X��9j���ڀ�
��ڃ�x����j��M�%���@�G�l��Ē�����š�B��(q=����E+FЏ���-(������ L
�G�w1v�%=K��bp�,�/�q#TZ��$MݏP�ZkO����\�����°�y���s?�)A�z�.�0"�r�J����/"�Q�Ëo����w,���pz�.�6m��2-Q$d�)*�X�h�K�zA���6�v�P�L*�Ø-N�h��HKT��a��3����n�����e���w�_�k�b���������|�>�ū���v�2k��V1@X�����}�����Y4]�5[��y�i��Y�U���Aj��% ^Go�c7�A~g�_�zТ�G!�� �|3��d�]�}��!�Y�����=� �`�7�w�~���[om�.����[�y���u�!>����)<�%K�7)��?=�h������92��]x8�s��]"�t"�M��
s����\�����^�h�62�lV���U�����f�z�Z��^:v�n��V;~���C������/����ܽ�$��PSe����3Ͼj[���ٕ��mo!3Yu?X��hwv��a���o�칗��o���$QUe���P�Ё� �Z`L�K;�[�E+!i��,��(��N��&d'�i���ܴ�,̺���f�Q�g����B2p��'c��PG����ͣCR��H�	1&a�<c��<d���|�U����Ӯ�|*~�\@� �#��U����e��C ���n�[u�, ���8;eS82�j���p�&�Uʸ0�L4'Q���
�@�����X��>�C6IN�����<�Y^���a0���xJ�SͤC������K`�(�QA`��l٩�P
D	��lY[1�:�c��B��T۵����T�(WS��j�W�j��[��}�PXŧw�:����?PlH��B�5��?T���V����N�(F=��}T���մ��=Jϡ�`m��4-��bZ�[ܗ��dȴ���~���0�����z��������hF	m+���䒞ۧ4�#���Ze�&�꼍j.$�����_Sj��}q ��u�a�`j�#�<���]FGx�CC8��ċ���@�`��y��7B)����;ua�޾�Y�B�6�}۬*}���L��S��έ٫��N�c�y<b��&�K`%@�p�wF?5��:R�z�|aދ@�eQ��^ڻ�e�
��d.�����|^��������.fl�Է�����`o�A#���E��FY킲5��݄ލ���k(�VպxܽH��Q�HGi�@����[� b�����/�k/��ý���� �J������*�jï��� �N�z�������/��C Zx�d4X�р��u��⑷_��~�m<Zx�([*Y�z���X#t��=��7l�AJ�sU��15J <�I#�,Yag���n����ОzyϞ~������k�H�x���lg���q� [R��H̠�3ϼ �^��n��^}�����߰����s���7����~ᔵ;=��v��b�>�}���n}��GQ7:}��@jt-Y���Y$'!���]�jZ�.��V�kwڶ?����w�=��Y{�̶�����g���m���߳��h��m���H�zU_ ����u�a�ٟ� �Y��n;��Y�<u�/��Ӗ�@h��}y!�X��g���s�m��։����k����ط�|�:���`�ӳ肔y�4�YN�-h��gc�5ȭx="���)2nd�d贪N�������K�B��,��d�d���5���ɐ�B.��j�w.��#�(C��I'�2��!��b ���WZ�!A� ���
�-�SS+�h�B��i�I�.�)Cȍy�L��UPy�b2�*���p��NN���O�wt ;�g��H� մ	5�&H_n�eNc4p&	�T��Gj$��8
�w�8�*�"�K�h�B_� �P��MRlm 
P�=��Da`��ѽ.���~Ň�
	�WsŚM-�뼽�m����@j%�P�jM�5קR���[5Y��Gs���q��δ��BWo�ݒ�Pf[�J!G�C����7wB@-���Z��Ԭ��>�U \���M�Ur�b���&œ	��p @���jz���6�T:��g�����Q��'�� �OR�Z��C�m�F�v�����CB���J9 �mo�FY��n��+�4J����j�����&4�R�� %�%�3u��0fՓ��ݩ�N�� �v�66נ1  ]�����j}�Z�*q*�;�R}�=���ֺ�K^r�'�!@(�x2o�D���a�I�r�� ����lxܣ��r>�*������{�2������K"���Бz�����fԪ-y������]Y7��L�SV�o�׿�}����"�	<���o���b����|%��/T�_}��x�m���������P�M�c��}�![�iQ�t�L�b,�n�ԟ%^V����.񠼻�Y�P�� �ve�ַ�o�e Kyxy�Q<J��u�9���<hss��)m{��g�>�y������k߲�뻤Il��3���h(zĖ/�>zi�����]݅�����!N2��������n՞x���?�����i��s_�����������������w>��נ*�;�rRCvҀ�4��f15�j4�+MJ��#�_����_������^ڲ-�J��
�E��7���سy�z�������k_�֟�W��}�;߳���W���?�������~˞�h���k/�r�^;u��ߧl}�e�,^�9��$�������~�1�Mh���}Þz�5����ǟx
>³�SŘ}�w[i
��_h@'"�ƻ8r쀍"��ކ�SM�O�0��󱧞�!uZ�+[��_��&u�^���y�c!+8{�`E�u��Z��w'��� �t`Ok�F�s-�����ğ�K�ղ�fJ�
��V��p�`���d���(�~���� ?<����u �Q˫��c�k �w�4�A}|Z�WK���|�G��WyAgj��@&���}@��L4ы���V��;�%U�:Z��V��i4��I�]���}�çM��Ղ(�Jsz5�B����+�����#��CC׻?|��w�����T��o��F�죏�YG�.�4a�sV�$m��Q��9z�{Z�L��H�O�љ����H-�`D������WD�-#	BqD�Byǽ��/�L�4�H��$��/lZM#��FP����}(@�� �h?�@�h�xRp�f1k#�&25�u�����)e�Ta8��J����X�Ӑ�PC�A��ͷM9 �:�}O�� �hCJ���@�_��ت��E�I(�!^����x�W���Τ�)���0~����*0E�M�P2Z�e���*'M����qq�0x�LHG+�w����^`�V�g;䡩�X����	m5�Q�]���L���e$�Z9�Q���+�R�A^+y����q���<��Զ�+(SF���[,gꁽ�WT�h��pH�3AA� #��V��٫AOꂺ�c��(��i�|�2�i�b	s�E��|��ko�������|�ТE�i�K�?��K��?��=���C�V��}w��j�_���V�����~���ڏ}�6[^�va�ti���+��/����O|�F�����fC���U�����sŒ �4�U;)hٮ;nZ��ǧ}�y�0c/�z�{��� ��vxeʊ���<���gӴ2��>jj�@�ԙKv��	_�OH�8F����C�i����v�]GmaN}�!���a_�����ʪ<�J�v�
Xz���왗_�k�E!�ڥJ������vݲSK�h9�rG&#Գ��䁫�M����l���{�[�����|���&�	;rx�>�����j�R~њ�{��W|)�ÇP��K�Tk?x�%{�����/�ngέ����|��v��'��~��O�cϼjS�+����}�;���X�"��_�7vϽ��'?���y�!k���cv��7Lk�&���t	��7��k�x��S�펛ݸO�i�q�Mv��
�LC�[�.�J���ҟ|�n��v���\����kϽ�a;������ ��8|�y��n//�E5 ���ȍ�+z��$ �FSY�#{����:r*�3{ L�݈��l� ��1���Aŧr��@�H�J�k��{�z�ՍZ<�p�wݑ����!�J+�y�J>q��FO� ;#@+�Qs�5@fss�"�b��z 2����2S%t̾?WK��iٍ�K�%���.�8);�ڲN�'�˵���w�>	D����5��K��i���Z0�)j���t�<?
d�; +�L#��ip��C5���A+�[@���^�e�x�k<^T���͆=��y��[���M�m��THT�O&W�݀�D��hh��i�<9����ݪR)�+�S^T�Y�MB�r���Մ	� a��J�]���fE����������Ccк ��N�~EK�7�� �O��(���ʝ��0�Ti!�/g�Y~w��(�x��6�4o�i��N6ɽ��p�՟�pE�+����x;a�d��0-�yD��t�b�O���Xïf�#n���w���仴8g�|�Rż%�~.c��)�͖,7]��ܬ��˖�rIs���z~�wʖ��W���Q"0_�
6E�ss|;on:a�e<��i��M�6��Ou"+��9���(C�; A�#��u<�4�`�Ҵ�/�jMUh�����Q	�� 
�y��]5�	 ��V���?���X!K��+�Ϟ�c�N�rܦ�D��L6�������ן�da���s8d��E�S��B��1�e�Y�E�R}�_�����o���l�4�&$�2W*؁C���K����%�P�R}e|x������W)���~���9��&�դ�>�2k�sx��.��hX�Ճ�v��Q<�B����3��~͊x��ԛF��G;�4k�3����-�x����r���ҡ�G������߽v����[n�����Ed�� `Đ��b(�	�P_��{��]:F\Gh ��a�n=�`��0k�za$J�U;zd֍����J��o<i��;_��E��;���iiy�>lw�}�����>����S�-����?�a��d�v���WO��6���w��o��4:@kB�>w�~�ӟ�O|�>;ybŎX����<y�W��uj�ڷ�|�{��I����VRu�A;3sE[]����X����ѷ^䛧��;ﱣ��)z�>���m���I/���F�4�.	?��{dZ�@K�i�+��?D�ERԱ �<�:t��b�@`O2xb�F�zA�Ǔ���T�o�e��G��'$7�Q^z�3�cP�J+�N���o4�Fȫ������۫T����7��`�9䴁���41�a��Z|�ԯ��d��ʖ�B"�NL�8��{�Z��J��:��i�!ҧ0:]@��PS�A������o���j�Ha?�̛-�#O��jED�4MǧD�OS)���������N�����V}z�<M�T���mދp�3(�y��T�3�	��(lKCU1r������!�P��,/��k�&�˕�@$=�(=�W�`11��}r�����4�N���1l@H54(lBo[<ѷB!ns ݕ�i����#v#�(�� �x�ز-^�M�]^��U�8�h�W�l~��yau��x���A��v!>�y��+ķ���-����36�:g�mve�3q h��9�✕1>e��4��㋶:_:���.ǲ��[MUK��<���y�rU8|����E����?�ds(�9����<y��Pͮ.�mfe�斕/�
��6�<(ܙe�E��]�~�P�/xSYy	C����,i]�\N�4�5n��ˎ[�OMŭ<�0������X�.^��%t�ߵ�6���w�y4ڮE��:�`j�3�9��	�w[x�u���b��Mq������Q�ۦ���j�$�E��k���'_�d�L\�]n�~��hse���>	�kէJs���_��^:e<�����޷ �%����������l��F���}��<�*� �m�4;?�ͬk=��מ'�Q0O���/Z":�;o9�C[�G�O�,��	$��k�'�};��'x�`G���Hs��I0@9����XդO< �+���'����;�X�L+��xN���Q�[�{��Sv
�J�5�HBWy�x��MY��'�^�B
�e�Z�y���[o: ��*��ӎ�5�O��i����oO>�<e�ٍ7���ב"
V��|�h<n�{u����_zo��}���U@�5{�� C`�Z�;v���u�<찝>���Գ{�Ö�2ʶ/x\*�� 0����lU���KW�s_x�vvz(X2	�*��,C9�j�C�Ĳ�1[���r�f_���>��������{�񙵶���^A��1�����IT#h;�8 M��5o5�G��ia_�Q�4r�ϫ]
4�,������Q����-�x'�Dc���+Eի:��դ�aJjmS=+����} �U�z-�������ѣ�2߫���1l(�k]�FZ]uQ��R�e�4zWe�w�Kӎ(ZZ,D�����"�/OM�C,�qa�|*��C5�O�B�4�g�x�j���.߻T}��ܨ�R]U����kr��b{�
��n#��� TC!?P��4`p/oqkcFZ&ڳ�}�^8�#}����_ٲ����f�nz����W^�
�:1+{���9���bf��}��bէ�H�x'��Q��=
�/Y���������枥�������2�{��IO�Q���=��gA�ځ���[P�Tf��j^l��S�=�/]		�bt*[ר<�$	�P��7���E9�r(�>qWY�59Z��TR�~p�G˽���P>� �ǩ{ԅ������'͡\M�&g<]�?!���ϓ7���H�(����q���Ky���gZ�@��Q�����Dd������B�H��kAR�6h) ?�����"Z��k���i���ݠɡ^��h`�o`ʥ�V�޳��=�,��[�8�"�MO���M�b��.��m^��@��r����K�(���Ks$^���1<��?i��/��7{h���~�* ���ؓO�d�.^BQ�l/�'?�q[Ę71������]Z۷Ǟz��Q���"|���H�@�QCv`����x�6{�����g��K�F�Z_�T�n���{�:k4�NjJ��J�R����羀�x�.ا>�A�ٟ����j��akc�8�=��k�r����_��?�E��#���݇7�@Q�-��v��}	��K��<��@Q�}r�00��r~^��5ae�zV�IrԴRf�<d~�v;����*�K���S���?}¾������ꇹﾻ����l�@�x��Z�^�}��g�_��(S*c���>;t�rܵ�?������N��"��q���}�CX���w��[P~�>c7�yz����d�����)�|�%����j��9kiRrbh'o=d?�Sw�{���T��gpζ��v��%uM�1��Q<�X�`Ͽv����!����u0H�0� |:�5P���j�nO&S*[M���C����u�1�SW��~�ZZp�x4�_s�0�D���#�S��6卅��f�^W�<�!FћFQ�>϶�oy�ey>����=��M��iY8�7�7J>��"��)�˂:���0�
v��Xqn��>�DS+���8����Ƶ�O�uQtP\�SF9�����`҆Ծ{�d���Nd�G-(]����TœR���X�mN>��&4���4[��Z5���Ko[���&���_}�ݻO���������>��ulnf�676QB�f������ I�:}ag-�,�Q3��ܬ�MUXYZ��gϹa���|��Q<\��>eeM��Cm�� �̺��f1vT^"�	�Q7T:t�� 	�c5Q��Qf������y���f�H��["��phVG$~ɿ��Ѽ�ɡ;~WDסD����oȰ�U�^R����P��/7�=�?0��^���o��,�SF���P*�X�C�
e�� nG��;x'V���=1O`����Ъ���SC+���9� ���M�L��0r���OyԷJ]kKj;�d,X[��D/o@���ph��\����۫/���/զ+�r@�(<2DQ-D�q:�m��Bz
��E��"�Z�`g-My�608��Z��P_� 5�,��m��s�)�N�}R)� �K�jjD��VG1��n<�)�*����Vg��=���FQ<�$�4
7e�槍bj`��=[Ļ�c��}Py +������E���S�|v:i�e�/�����h��s�4;��ʃ���gN�������^�y��l��ܪ�ٹ9�����]�F�%Jx@�xFM����jJz=�O������u�Ze�2^�;�d7�xطv�Ru���]�~���~�MO/�Af�IM��o8q�Z�t>�%�ⶳ_�s�ϘH@�B	#���\�
%�	�Ӥ+�L�k+� ���ju��]��ڴ�� ք��w�8?��u5o���5{�ų6L�h�M��7��b�SE�vئL�@��R~�t¶�vޖ�3�e�j�L�v�����]:���ޜ#��xR �3��ڴ0�W���ѝm�u��@{]��l�1R_��C�<y��Ƽ�d�ۼ��	!_P:��i�����m��%e� G��!KNS�vw���U�K�"�E^�Z83����5�߾ߩ��<����(�qT�pT�Ľ�qE]����T�0��}5���l%�gjm4G�,�M;��n�r	k���Eo)]#��.ը�,�E9w���F���y�(J���cS��V�݇�<Iy��h�Fv��oP.��oZwT@�@�Yr=#����d:����~�{����Q<�/��ϟ���-],������pCS�j��5�P�mwg4Y"� �,�u���mnvf����7�ĬV@�cM!М4�b|��U{HJ�6g'��[n:l�M��y%m��>5*&L$`=В�s����|4@���
��F_�"M��Z�0#��p���Ȩ(m7?�z��}>RFa�R�c���LB.��!������Mt�$n<ha��T�/��v��>�r{(E�3W8�WY��y�1g��Ѯ�ԇ�C}���=-�{:k���ھ5�Gg���w��ҒDʇ�wi��v'���c�Բ5��BT�Q"���k%�Ђ��.�W;)� ��ig?؂����f!�et"�G�A���]|�5��[�ẋPa@��ZfJSZ4��#�ZR,�"�D�Gڒ(���K܎�D7�Y��S�XU�fu<�n8�����s��|�~���f���\�8�q����Ee�d���'��fY����j)�������.Jq���Յ�! �"#�hx.c�=U�pjʮlaX-k�;m��&�����N�/�d)P�g>�Q[Vs�tٴX��J}�����^�H|ӾRC�@�Q$Ä�m���z�V�s�� ����F�F����\!~�,L}C~��	���'�Q:_�9��{{��%������S������-���-��2�N�K݄�ɹ�[���6��v�J�jm5�M��x�t��u�.�Bk<A�%K����J���s��;��"F5
0�4��^9���i��u;����M{鵳���g��>��`�����h2�M�]�,Ʃ�4qj
Ǵ����?p����S�><�~
�efX"?c�K|��g�h�dpE� �B:e+�nZ��>���ͺҍ�xĖ������08ڥ^{�iq-%��`G�X�~�<�0Ț��/fHy�p<J�� �Ш���%��ZZ�S� 
F�H�p04�R{j��V}�*[mԬ��=K�Ect ����ed�M�"��`9��hʏvb_^��r>�Q�h]�7���3�idT{-f��Uk�뻕}��	��Sח�?���w�.`��g�!�gy�b073K�'����3�H�s�<Ƶ������nź����9�e�0�w>��إ,��
��K6�U#3���I��?��Z4Z���T)W�=��Z;Mm��O+2����GRg���j�����Z =-E1� ��z&�vDe�������5�C� ̵=<0\[�QW��յ��y͢p5BP���J�ėR��())^�5�P
���R2p#�K�Y#W]k4����F�ʈ�?���T�H#���<-!�E�5����<����qкn�%���8y�{a��Ⱥ1�Ss@��Z~@�B������s��V���� � �~N��<D�K�F0�گ+T?A�R��π2�:dĵG���;�<C�C=�Q��#��r��X��mg�?a���>=�HKڤ���������lCK�ﮭi�-��"�9A��ViG\Q�xX#l3j�A��T�{���M*]���'B�]*�F�;QYl��ik��i��2VfFںH���c�46Ϸ�6J�^t٪ݢ5y�Q��ܢ��Ї�c�F(�����m5͕yń�%2V�V��~�D�l�C�b����ڜ����"�m�^��hu�� i�^
�MYbj�Cnz��HZ9U����y���]��fmo���Fĺ���O\��ao?�d�!�%��[� �f�����9 -(��F�$��� k��DK�
��.�E��Z�|�¹��W-9uz�ؖƏH'���פ4ѿϳt���TM7(Z;�xӶߍA�(��֢.���U�������&��,u�������j�������
K�ϢH��:14�f�,��8��������X,����a`0Ez�.
D#�Gx#�X����uh�7AiA�>��OJ��4�ϱ�E_�M�5P*.C��k���s,[ ����.��ĸ��cjx���L�5� j�%�^�ɓ�6�ź�b)k��~ՂC|	MC�)�mWdd��f-�`��=M����gį�2����%y���B�j��(��s>y\�����Ps��E $�0õs���<����tÏ�c���j��8h5MEy[,罌ihvlu֦�)�6`���R}�A(�l֦�v���� ��y���.̖�Gtj4X�W��Բ�E�T�`Q~EІd����8x�j�~��J����Z�B�9���Z��q�cɖm�n[�JŖx��q�W��mno{{�K�$@y�Z�R����.��*��Ȝ&	
�K!�'��V�u�����C�Au������!�F��\n\Ԇ�ByB�w5�͒jf��g�+d��난<�s�֡����<q�zd�Իr����x�}�V�=pO��q�]a���q]<ϓ2������ ���-���P�r�u&�ބ�!p]��\Y4�JfL�F��,�_h���G�`fu���5E���4�AH}�w8��G�&�C���C��R�[�rH�-���`��05cC���v[�M��>��A凗�!;��[)No�|��9�	�<����X0�
�T�����{̠��
(VղE�,X��{��5r|��2�<��Fx�C�_9fg~�����wN�ړ�*�}������b�[/=K�0��9��<��8g�{������9�ے(}m���v-��h]�בT��q�F5yiq��C,�"#�l�5�/c4��`/y�l	uB���*`��<�����7-�Ս�@�=@�^�A�߷�kE 3�-jf�M�w��>^[o����)8'nD�{E�S�V4 gp"�;��Wk�<r��4�m���A����Cq�;@8zP�D�R�ꊨ4���-�,��u)��fg5�K��q���EߵB�5�W?�qi:��=�;�X3�$p@ԯ���jU�zK�ZL�S�E�%�嫑�z_���R�d��T�;2��C����HK��ˈh����-�T�]-oEM�����l��[�V�EJ�R�F�Fr
0hzS�<��$�}��W׈!"�D�,<��#뢽k]�k���6J/��LL]3W�u��q��S3=����Ϥ�"�o��Gu_�<N]���/�f��0;��50E#5�����H���q�����4�F;�k:��i��д��C5��?Om�%��)�Z��R��^��yu��1*R}B2r!���L�%�=�(MXV����к}Y{)�1�8�꽂^�ٕ����Ǎ�d��q\��=��oT�'�-�!p�Wς[W���=�M$��t��'�\=�3�?HW�|�[�p���'�R�gI����92>]{��yx�)x�q.u��D<Q���T����m��%����^���Pߪ�$��y<�YJIg��ԏ�7�~�z��]�̈́������e��+>��`x�~��1�/�<�З�7C҆\��|_�>
2��������������84|Ҵ�r�I���>���},K���F�ɸc,��M{��}멷챧��7�8cO�p���ɓ��82�r�Ɓ��Sa�<��q�����R�AY��~�<�u���k0�}��k�݁�@>���_g��Xp&�A�z�I#�S��!��G��T`Pcx�n�ya���P��M@􃑦����yh/��� ^B�8�8 ͔-S��T�`�z�* �|��|��V3����>:Kv&��+mh~٦�O��'���7�vN��i7�m��TiUճd�iP�����5M�Q3<�����U�_j���ˬhoBt���$x�)�Q|���%���ߝ�I�(]��2޺��+m����"�Qcb�_�m��X�R�������2S�4|uec��^�UHdJ��AP?�~�Rr�V�U|�ҥ�"2`,��IFϟ=�N�#H�aW4���K���YGFz4��좟��R��1mB�������S�Ak6���Ռ�M�5�o(�(� ��5u�%Sތm\��FN�Ѩ�G�� ��9@+�soS)��F����+6�%7�o��Gy��X�S�|Z������p��R�cRL��ܨW��e�o�J��S��*V��K�j�<=Y|5�i�(L���bw즛��B���˩&;����$��4�u��7�fQ
�q��(0��Y���]�ֿy/�͡W<������s���e��/�����
�g��0�C%H��=u�q{:2m�\+O���|y~����iN��`��� @����虚8�ί�;5�����)����8�?󒿧?A�q�9ȯ���5��Zg�v.�7 ��	6ǔA����+��q�%-��G`��X����T_��o�):4�f$�sbxE��ƙ��7?�=g��q��A���a�>iV�������3�ϙ��Z�����S&�*��^���;�U�*�ЛQc��m��+�k����=bu5���^A��qU������}�)�	�Ys������=	r~T6�+����U72��/�C�r+��yB(:��`3T}/C�|c Fc`��A}�ʞ�||4���V�b2$��v4�g�!�9fN�-L�C���h�ؠ��Ȩ}s���A�h�Tߠ'����}�u4�	�'�7eX�C�_t �]��VNJȓ�a�P_�{McV�i*H͏x�{E�w���e��B��淉Κ��Vw@�?4Л��&z��Eh��T��9vxM��v!ה,��yGM�jf]���Z<3÷)��t9"o��.ޔa�P�Y`������˨Z)(�/�FY��FhÞV�����0z��H^�� �fD��Eʫ�yͽS���~ ����%�&ۄ�.hS�����j�5QjZ���9`A/��l�t�&���i�ܢ�����L���=x����H���Ϳ��!H!{�Ҿ=�
/1c�Ҭ]�p�3%�NꪏQC��(����:��H%1��~F���R;�K"�[+�h~V�I#pZFGC��߄��ɛ��bκ���H���)�T� 4&����:����%���7�{t�QMj��*'���:&���?��R�4�{T�1�c<�"�C����m�{�C�A^�֙8�#�=Q�Ϸ�F`h5�^�7tׇ�sW�j���G�{:_�o.��;O{R��,�z3t�3�ͧ�+j^���+�)H[�ϡk�<�����Jςp��&t	~eA���Y[(�k��m�M�.P�B�xlxZ�B�%L��� q&��FCς��9 � ���?�I�'��4m��L�B���&\3�JC%�|��1kP�?s���N���S||�r�1
�>c�PC�ēE�DF����E�Q�Ȏ��8�$���x9y=s-�a� @(/�C��A[�?�"��M�dp4��7�������A��/��q<�-� ��p5�	k��`�{
��Px����M��H������Ԭ�7��ZK	��P����:�\�r�( z֦�i۹|�vȅ@��\��T�E���N8�򑓒7u�d�xyR'z��W�Ҕ4�g˔5�"O`Ġ
[ۨ�iPkǠm���'}�R]ս�=-���V���y���-o������xZ2�<!w�' Tk�By�"��CuS>|�G��e |Tx$c��4�)�����U5L�j��4E��]k ��U��Z�$��{�y"�C�p`��0���@�^׊�����O^�"���8�C���ꞃ*�+L�g�U�ҹy�w���W��"��M^4PM�td�yV�Ļr�����p��t~��[\�u��=6x�P�wԟ��'�o��GU��~���=��K�,]��K�0��HLOK���(D
F��	�CW#&���|�IJ�v[5_����6���0f2�0���^�[���3
��mۈW���^�w�pO!��`ʱG���婂�٥[�'��;>zGP:T��9L���w��R˓鷚Ye"c��y� ����������/���oģ��s0T�z�4 t�������J@����"��on�)*���L�U0��Az̝̕��w�����xA�Hg}+C��
H3��v$��:(�ӆ<ʘ;�<� ��Fu�W<�ɸI؟�1���ƇzJ�j��O������� Q5��Q��W�w�Q�B�^W���:B��`p����)�>�T��Gj�!�
�ꙿt�����u���x=n����$?�G(�G*8�����q�y]���Q$D����A�"V��~�p5L�GI��8�乻vGx�y@��x���G��8]�,ޫ�	T���A��!(}�XɀjRM�jI	�)5��?}�G���*\�"σ��&9T�`r��uK��кi���zfcȽA�Z��o����c����[ �]붫�Tצ2=��vEZtk.�<<�����x�{����B�G֠�!�j^�^W�G���=0�����1��ӰV��xC7jX��dQ�
����֑A�-i+2ţA,	h�o�ټ������"�j�OO}g���`���SO�
k���A��eEW�ӫ�KLC-��qDqF\ �MJ_{w��{�� ��/��x�~��v�!-��zՅ���5h�A0|LZO�&��S 3�"Kʳ�~R����g��������9ik���<Bo��t�{�cŇ�T���RVr�4c@e҂�-�Va��6;]��n�{��6�����K�B`����ø�vv۾��Y��˖g�����&<b*C�LMMa���$��)⑼?2�&)��-..��ֈL���x��H%�6=7��ݳ&�|Í�me����qI�E���~ס�ֵ������~w`�;U����Óн�<P�� {�L���F�I����_�ko�&��U��F��B:�`|}}-��NyMs�F5��WHW��C1�5Γ�%~)%!)n�&�k)R�tR����_|�+|EԌ���)5&�4d`,����ޤ�{�@e��+>���^�����
��P�7���6QB���7��r��;��o��էc&r���H$VBP� &?�ʠ0���r��?�^���������w�k�f\K����L^�}5Ny�J��=/?����?����:���鏌�����k��3�4_A�uL�*�Sp���}:_���Ư;�����del\� ����;�� ~8�q�U)u��W0RU�ε�E����۽7,������$��\�-���|��e�>t�	��Č-N����l6d��);�������e��H�
�����,my����u��綣�TNYtP���E/�l:�幬$�[o\�G�0 �a޲��(�
��D�ֻٱl�]۱*�b�^7�tc�ԈƂ�2�TmЬƬ���F47Y�i��Z�۰~���a1j��<J�b��n��Q����ѷ2��
�Ӫlڨ#��Ĉ����֮3y�Ƿn��5�i׌�vL��8�Q�e9�6���ma�0�}��@���-��>������\X���h��N�����u��o�L���"oN�6�n�I�[��W�(�G���׶Y�{�i�6Εl��VSzڈ@�/M�2ٔ��N�ylG}x�S���n��V ӭ�ʨ����'�K��i�������c'���_�uE�Ǡ�Zm2��e�J߮�_A�ðx"=\P\���}��	;u�-_xZR���S�$��w��W.�Ze�~�g?b��1�O&Ө ��!���A�%ø�0��&6�b�g�;V՜+��:Ze(�7���'G�ß��X19!�����L�A���c��������;��B�BJ���d�.t��TL�猨���ր!y^���Kѽϔ����DPyjˣ�(HG��kb�&t�fH)`���>�;( ��tKC��q��=��ȇ��)XwRRY���U���I*͓�CJr`�����N�f�;���Xe����[�Y�Z8Q�>����@�F�S��{ޕ2g�i����}�~
ٯ��=���;ݼ�����8����u�������J��|(x���\w�p5zq|y}"��	���x���t���G�C��������P��c��;ix���>O>QyS<S:��i��c���[O�1D	�/$� ߣ�0��j��HB�T��q�|�o�#~���
M�j��Ye_��S=h?5)pT�O5� ��[�"I.�\��@�4��������ɋ\���?kg7�����2KV��,���!�8��m]Z�W�mz�����詨<�`�Oەso-`���� u /�}'��h��So�c4�Ƭ4�`q<0ͳ���w�w��W�Q��1�f�V^\��F��ق͖K��+�ڰQE'�+RE�M/�v��p�[N�3o�l��ϣ��(������^��M�;��o����!��%�S�Η��K�"�n�μ���7�&_��_�(�/���]|�u�a�Ղ�d�<?�}�jqY�54�|�y ���e8<���]\�Éi�ڕ4-!�.XpP��.�J����҅��()���Q����[n��z��x��Z}�P�~���j?��iiJ؈ ��¤���T�3��3�lD���C�`���1���������e���D���.K�"�f?H��V�I�c�
�{W�$�d���¸,�<��+��>�)���^�j��YIE�'���x)ʔT����a�y�[ln[��i����m?�����m��_��'9?��m=�=k�4���V�n�<��F�� =i�`7l�8�\�
)�������>����w:L�?|���+-'��(c7I�j�?����=���;'��e!�k�כ��k$�F�q�f�G��ě��3�)�Q�룝b#��8DA�
�![���$h����������� �k��Օ�⾂�)� -=�*��!�G���q�I(���T�"B���d'*# ��\+�E�g
�-�A@r4�Ã���ASX�����Ă�X��3)I�jT#��y}������� H_:C�=}  ��=5�լ}��E{�E;^�Y���x�+�5��Bvl*fɾ��=ˡ���a15�x�w,g����0���<������������u,	���6�][*�����e��@���v�г���V��-�7N�C7��O<|�>��m6[Bj�-�0��R.mG��M�Hg�џz�pa�I��v<�h��ֳt4�w.�I��v`q�7Fռ����V����Q������L9�'���"���TϫJ�ڠ���x�Z��_��VLS�x��^�����>�/�Y��S  m${hq�槵�I>Q_\�ԓ�9B�a�2,�OS�]��j��(��-!�b>g�+K������UV$�� �Uː�C�mv6�s�ᙇ4�c�ya�H�Ð��Z�M�*�3���L*��\�u�h�cZ����R���sh�C_r��}�����,�f��^���-�|��S�~��"t�ϻ�Nӧ"h�H������T������'x�%l4[?I�Ա����2�\���QsD&G 6?|��;��p4�����;��� Bc-��I�h絁"ƭs�m�
�{���W>o/��߱W���퍯�����/عo|�.־�v��_�p��^����[������γ߱:�l��o3{�0=Sɠ$%<���N55�\��2��ϋL�2bA�UvD_ �7	~r�0���`~�Uz뾿3>��:��$y���f�c�T$��� O���(�;���!	D�s\���o�c��y|�%�"v-D������Ϛ������[B�������P�t�$��ɏB�C�]������C��$&����8(�q\I�	A�E��8�����B:٠A��9ķ!��?=s?����A��Ǎ�?W߲�'�����7�����BݡH�y�k,�3ܫ�/Y��@�2(�)<����w����X
�)dA�q	�Zyڔ���GO��h˙ 7�?p��,zH!���&��D-���$��<��0�y�-CP~����D&�w׊�0B�:z��=�ū�@>������u�L����b�A�-�����;M7h�~\#���{2�'����{��D�s��D��	jҔmצe�x`ޯUj|^z7�����䤨�N���2:w�]�ޱVì�BoN�]�_�G�8�;��CF^�Gs�Pv��.GڷS BN�G�������x�}x��i�L�
�����@��RPc2���k��OG#���Qg��Ts(�̤���������M��Y��X��u��#����>�F��z�^zk�N_�� ���Դ7YjR~��)Tu$���ry�?��h���q=e��/��2Z�K��h್|��l%4�-kS8�e/��#���*J�2��@D��Vc��~�����7��ם2rLvU^ 7���kW'ih�t���1�B_�ے �P�E�7�i��o�n�_~��=��m���UϽb�3�Yw�,�Y�xk��Kuw1�5%�޷hSk��Y��k��5ۻ��m�~ծ�����3)�����ݶ<a������m�|��>?������6��<�Tؒi�d�ѩG����*�G��(�P��������6�ղB�w��4r�xq?|�S�g���<*�8�M`N�Y!�<s�.lR�pYO���<�ԩB��cxK֩��ԇQEXk�PGQ4`x�[�O�KҠ*��yMD��6��;B�� ie
W�(\=�w�@��#�w�׽ x���6#�M��a�] @�
�]
SA["��<;���IEhp����j����2�d���)�+��dSr�����itϯ1D2d�4�ݵ�eRd��56n���(���my�7�OZ��C�]��nH��k��8(����{v/�Wm&�<��bߧ�{Cx%�<j}��2Ӽ1�����j�:���t�6���l�����~�5�.X ���KF�� �=E<�C!�0h�B��_��+��o�b���%gME>���\ζ66l{{�lA�HҪ}�S�P,��҆���#m-���z�����[\�E>��6܀i�zT{Ib|��1U���bv��$�(�����7j��4����.[ew��c��t"��QUW��ꪏ8�x�����Z:k���D�:�07}v�ԛ>�@:T]ZvO��n8~��*|�,< ] c�G���~M-?������%�<W��Av�)�+J>�us{�|C��9����gL��no�x����%dmxeJ;c䊶qe�ꕪ/����z�[+�L�,�j9k���-�BM{��#�Z�W����I������_{�~���(Ȗn��~��C� Z3MS\ia�4��T�T("uz��r���IL�xb���d�5��1�;�����>���u;X����?t(��!~��lP8���@�s�=��׳��|^9��G�jF��Rľ�+y��[H�E�e��a�L�Xo�=c�����3֮m�yZzG:�VR(���$2���Ea��<�:�z�d�a˚+��U�.H�0c��V>p�򋫖\:d�Lښ(	m������Fb��"�?u��ƉS��E�#���=xh�B���̅�:�e���� )7���b����Z�2y��*�vp��@�O�VF�Hz�>��%+'�����:72C]��IHIC�(<	I	kˠ*B��t�1���GPǓg�'{�W�0�[�4���>��ߛ��q�������A|�4\����i�ޙ�U5�TY$=�ޙ�������~�o��kG��J��q͵;y�J.^���I�&�ݹV��ϧ��,����d�H���>}��g���D�!��ܪ���^�ͭ=��擦uռ/���ۧ���sĬm�ⶴ�`sss>�n�ʺ�c<�mY�^�����E;t`ղy�H�e[(ޚ��)[X��,��=� Щ�W3���� %U�᷿������?�H�nt��6��/�ҙ������OX�+a�X#��r`�m���se,��E�S��j��⼵Q���/���R�lC�����hz~�R���yp	�Z1h��L�n�29�-O���_E�Sǘ��Kh�A��G�<7c�W�l��y�Lx��$Ά�c�5���uԱ�o�F���i�k_�:����%)g�x�ܣ��[�8�t�vk�?�S96.��ZuÍlX�Hc 
JfZ���F�bW.]��%_I�D}x19x���Fu���!�0���Y������ԽV�Ҏ/�Ei����Y�ѰW_xÊ��Lx��Ư��� ����;�駟E٣�x���	2�UD4�R�M�T��Z��w�#�Q�PM�7YIp��mKc��vA����>���/DEv-	�����.!����55��Z���9���G�������˯�d�(�L�����1�=V/_���_��/�`m^���E;��^[��#�J#�P��?Q?����d� z����D	�P�ߝ``�;BG����m��{-�z�b��F@(�v���	�N
��E�Z�2~x����y�{k�E�H�ʳ�oZ�c��<y�u����O�d}��(�z�2�+�ɇ�,=j�?����K�)�n��:�S����u��E-�>Tn�Mpȋ�h�8���*�+�2\5x�3x70 
�D�������x��w�e�*���+��Cu����x�Ұ~ä��������ם^r|�09�[�<�<������u世O_=D�^{W}����Ǥl�g� ��ɔ��f���?�1�s����R���<:���u����b�?��u��xU�iW�k�����|`���~��6].����U���^#3��Ҳ��)������a�����9}��(^�|)/�@�xy(֮ {�~���������3�o� ͯ<{�~�|��[�Z�V��S�V���N��+�N(W�I�H�7�u��TkD�:�ZP��l�ơ�Z�(��0��)�С�;�"��C��p��-e����6��'T�u�5��UٱBJẾ�����3�&=��N�R�%�ء��Z+6�e����f����u� ��;)�!�Q�chK��51�����T�SsV�b�ЬP*@�+���x�4�^#��'Z{Y��j��v�Т�	���dԽ��/�K��Dͬ!���őqʐN�x��\;�I��A_������7�n�d�B{���2E>�w�����X�D��7���[ ��M�-�e,���&��S����P���%V�c�U��S8��:��)"MX�yUT�)
�}�zm;xh��Σt� �C�A���q�`��Z��L�z�<�����4O͙6���C�Bv]?�&��6�X9��U�=�^8m����]|�{f[�n�2�,���ī���u���M5As���zsHI�h;(�l�	��+1���k��6��c9eh�Q(٩[sw��7�Xm׍�VW/gs &�� z��D3]ԑ�} ������&��	<�{}�(���FXI�i�s}�^����J�k�3�)��]�s�"��PH��)gE׵���Gؾ��� '@ ����NiS�~�F]����#����������挃�e�5�XMS��|\���*!hZM��=P���E}s}x�{���+� 9�u����Ǡ��o��h����T����ĕ �Z@C���͛�@��Y�)��Ix�NC���C����д݋Z$b��=�7�3����FgO~O�/Ϯ�k��͓ދ��'y�澩p����w�*u+��z3<�5�g��_y�Ywi�u���l�N�t�>������n8q�r٤>�bw�v���[Y]�#��m��l��~��|�	[^Z�F�`����.�I�m������];{��Rq�wҥ�0���V�����5�Z��45H~����M���1�B��O���N�)^衈5B{AJ7���9���#�Ac"�b����h���7��먉X�X�3 �P�wԽ�'HJ5?Z���2p�y�@��%���8 �2�!�k �-4"z8�S>�vL����J�����Q����+��a���Py�?��F��'�MzS��Ii)4��r� @�)r�%)��a�VZQ_��WQG�0�,r��B�h�Q�ڸ�<S�:�����5�}4i�%����Q�����K��1x�n�J���/�z�6�'��5�N�������T��V���V6��Z(�f�r��Z�G�,;d�*kBc�J�ƚ,���#GVa�ޡb��/$�������zr�zM�������,�Wq�'D��AI�� �J��������s4�%�@�_�h��{�6��������70v]+�%���Qt$w�#� �Rj�WǮ�D}�,�ֵ��D�J��DQJ�~RM�L�M�{R��Fe���;Ͷ���$��0��
��x�����Dk�	�x�y�ᆊt��΃�/���f��^.|������c�M?9�ݤ>t\�3��W��i����Rq�A�n:Z ����uu�1�N
Q\�oW�62vB�E�z�_�]��*���q���Z7�y�3����%1&^��׾{g�'�*��o�y��t�ߓ��@�Ԕ����;�a�z�*�~�6�O�� �Ƀ�#C:�/�J$�N�� �ڌ3Jл���k=�kԐ�O<!�ş>�S��A��<���һz��(��Q$���PQg�߰{N���:B�����������/~�x�!�ۣ��g�<t��sϭxpI�?��P�!2x��i��m�Q��h�\!�D�����*�����63[�3<i3��v�=wۧ>�)���>�2�����lzz���=�=�:$om�ؗ�����%����(�F�ʊ51���-�(��J�p5/P�1� !d]�D�+�.ߡ#���Eߪ�L2�n"�5[�E<�A��}^��'�E�!q�b ���{5�M�w;����	؋��r'��;Ǡ�o�t��
�KW����7���q�֟.���^6����C�92"��!�V�V��ĭ C�%����g�O�fh���H��79�k��ye� f�SMS�Sք>��n�����{ځiɥ*QT�e�E娑�=
��	�{w(��\����@GW�.���.��F!KMA
����"Q��b\���iԦ<����IЀ$�DD���K�r8�u���z��CsY��u�^B�@٨|z��]]mE1*M����Zc��ڨ�1��gc=����ǿj���i��oY��gS9<�x�Z}ͯѶ����x�1IТլ�0���M�,���`d)�$�K�FzM�s���e�,�fS�O��UJ�,����dO��+Vy�	���?�ƫ�Z	���ԑQ0`B{t����s��R�OPt	��8�����<�u/����:�����\n(�A���(��Mx��8�ad��jI�����2jJ�D�>F�-:�	k��m�£�/����G$�äUu����=�c���R�Or�"���P% ��oy���1x6
/Ed	�_"-��@��=�=���4�^�>��j�#x��D8��j �C�8����M�h�Є��d��)ūe�nl�t�|ۄM��$}���
=��� t�]Ak76�O�7<hk����r�{!��C��w�~��[(�&2��@^��tjS�6Z@�.mbWA4%O�3������ǒg� Ң�j�S���(]UyC�Rma�6]�q�:�:��no����e+1fŜm���+����z��r��\�lg��P[�h4!r���aO=�={�����U����]n�=d�����Q�:^z�E7\��'�����T�d3Kn�J�M�[!��KӖխ�s�{oY�vΊq(�ٷ�|�ͫ+���w֭�~��Æ�s��Z���<�~چ�m�~��r�)���r�q$z�]uv/ۨ�m���1��J�B��0�7j��P�	���B)iI �P��%�M���*_c���m�o77mT�6��[��U�#�7����T�����ٻH�X��eٺ^pN��e�5��/���x��x�]o�`]��A'���9�P�z���2�w���l���b#X۲^{���l�Z,E9c��M��r]ڲA�f�v�Rj"�@1��|h��$�S:FΚ����J�%��������4�@#�H]���*x��eAh�
����Eґ�ʓ[�^B�IM����Bx�(����I�����X���1֓?t���/}���iY�D�OW�BK:(�#w����d�l�V��R*j��[{��x��^�T�Ra���À�����' q_��&)�l.m�|!U����D�b��-�2;�R��N�[n>l�b ��0n�p�DiA�B�#�QMqB���\�K^6���kv�Ǭ��6�|6E�@E��+UǸ�^'dL4o�i-:����1����Q�8�_c7er=����-�+$	�*e�V�@�j�ˣ@��w����6���F������A�p
0��I�Z YK�i����0�BY�Z�W����Bδ	�PAׄa4��:v]�����ߍH+4>+(m���ڍ�ЏM�]+rDQ�J�o��=pO�&�B;��(�8��_BA�Ў�P�]��ӻ���x����`=-��{�iC[~�	=�� �Y�gJ�V��ﻼ{}蓮�A\�k���%�N��SS6 �q��4F�)�/Oa8�JI��rA�A,c!�mF*m����4��5����X4f�����:������}��O�믽�{���_����׉��vh��-O��ޙ�Z�Z{��W����:�[W�6=�yas�m�[�ff��S���R���_��.ɉFc�ϩF��F�1J��3�'�aHU�l�e�^|�͍��	Sxq�.Fnбd���X����3y_W6�'[��M+���p��}O6m�
�(z��,6�X)ݷ��Y���;;�m��jVƚ����h��4 �Ҕ�ޮE�yp��=8Gي(��_�-��ќE����6e��%ou����-�nZ#!�l*dG����%F{��rnX:d�}q�A��t_��c�ac��M��b�n� ��A�X�G�y|�4Js�����,�����U#���\-z?h�V�u�Y�%C]7�>
v����P�N�*S�s�
�2rm��۵FלC�S���Ĩ(�F��ʒ�*ћW�}L_��k�����+�gx�;P����a;�8��W����!e�mA¸u2��x�yac6 }�z�۶��s��<���'���pg�h�E"��2d��+Ĝ�)?�tsv`i�>���3����������O�����g���_����G�;����3v�P	䒧B1� ��<D*\�c�+��s&���{�������ӏ[��Y��C�F��ԑ&�^*gД;>�)�
l��1�~� ���=��.͏����ש�������҈�t*idہGL)\ȬӰns�|]C����4JH[��P�!�BXg�~�z�(�(�<�(�Y	����E���&�^&u��!]��)q�{���P�>x�e�6�c7�����.3	��>x�����|�~�4�6D\��E
e�f,Z��pa���9¬ErA�r�^4?c�Og��ߔ#(���ĩ<(��\����ޝ�a�k�	�u��K05C��x?����p��%硛�=O�C��ߜ�I���^���$��R��k7k��T��桉���P���XA����x��"5�y睾��ɛO��Cډn�������Av�v��q;pࠝ;w��x0��yW���|Pm(�w���"�0������t��"��B��㌢ƈ���WZ@��(n���˦����e2� ��b�b�.���� #��g��ċ��%�ˡ����0�8 9�P����[�( o�vq,ܶl��o4u*Oy��l�Q�n���ڤ���nC�!�v��[�c�FK\FT;�9@Ts�	�@�[��ڥ �����t�4MN�'C�Z5�b��I76�^l�\�Xo���XCu���uM����Nj샔�0��D�D��^���>$�re=�k���Q��v5;�fZ�sT��P`?<�>С��ɩ�F�p��A1B:�ᣝ(��}O&MtT_�:ڵ����8�~�0��gW������/z.�?���rUR�:�3%E(զ�e�m
��V�������� e�ʃeG
Z�� ����F����2x�w��=�'����,ZߵY*7�K�w|`�T4��|�#��V�٬�  ���A�����o���������/ٽw�j�eޡ�{-����.-�mn6a�l������ D0��8����Һ'�Y�ET�r�{��_����V��2B3^��20*��s*(��)����
����� �+�������˱rVI�����j�sv����8`c��$�����1c`��`�`H�Ƕ�9'�ԭ�J*U�/����k�[O�n�����tt������}���nu˟�YtI�����w���-���ƪ�+�ڕ�`�ޣɤZ��<��&'.����)gQ��Daa��&��jJ��]��ZMA`�Ч��+�!K�Z��$h]<��dfu��l%-'��NTr�W#sY�9YyJX-��fr�(�ZM7A�#�ν���d;���
|uM�gZ
�z���$�g����>��D^�P:�vR��P�"�K,��T���;uˏ��oT�H��_3��b �����3�)��g������u���ǼO�E`�r�]S��^r7�7-���|�z����e�,)_j;'ՙ?��Pc�NOk[ŲƜEX�V����Je���(:���a��}�]����b`��I�h�ƍشi:|���,�Q����_T���ކ�k�b��Mh# Z�q
WM]�ר��/�@�`!�շ��F�L�33�x��\V�dM�m&+M(Th�iq�*m���[PV�j��&�W����;XS�*�NfP!C�h���}JZ�~�|'�ټ H��Hrȳ�R�<_aÖ�A����Ūx��-����-��a���d�UJds*S.ЖB��RXx(��g�qU����L� ��ڍ�#i�K|?�$���QaѪ��[yv���w&�:\b��K�#�;�8ϕ��|��`-2PJ���Rf�[�$u0V�lG�8��H�ժb��P�fXμ�h�!�Hi1��h�W�TW���L�Q��8�uuʍU���4X��$���9��Jh�Z�Bdhs�喧6�g�]m\��M�_��j,��AO�h�ѧe�ɗ"0h|Qy�om,//�b^Vna~g�z��<Wf-����*�m�����C¥�"K��2ISTR����`]X�zv�܂�o:���C������.��o����/����������5�E��D�
��ch���^b��T9�h _���	�%�}d��"��ɧ�@nb��^�Z`��U�J��Gm�u�A�^�__��z�����{y�����8�RKHi%dE���Y@*1O���]L�\)�I���W����!�Ԕ�	-D��*N�� *ML��}ur�85;Ik�՚�WR��?%�׼����k�.�]Y�FYq�&U�թ�f2�Ge������H�Dba��z#Q˕�_%ݙ��T]N5%������(m$-�eb��M
*
�
�o���%W�Wuk�V�SI��X.KV/����XR���e[!@U� 8{1�˞0��U;�o&���T>�^��U��z	�ZύI����VPZq[����-&-`�T�u*-?&�;��<h�Dޔ��Ũ��'y�z�L��l�.�R`�	��	��Z�(ޯѦ��sʹe9�ɮ� �Md�Ů�y
c�cM����9L�g����%�7�+�h�j>0͸ɹ,fH�T�� ��'��f�Ia>��IZw����� �{��\a$�U,�ʴh|���J��(��u��s�
�f�SU/��>棝�@2SG:�b��	�Y$�*Q-lw� �Aa�Ǽ�qy:��yZ�Tp����ոk~ɏ�O$�XdsKl?Z\�urF��C��7NOO�z<�x�6��Z�V�ó���y�J���ׄTf���h<�R�X�:�*[�#��O����3��0���QbPm^�Cr�\�q~9�[Y�Bm�H��D&�x���Fdxi�^yQ�3�mU3�D��9�4�S�
�E!��s>iL���"gS�׳��J��W��c��h256�gs���^9�䥱5�*O:������	S�����`��ax�=��h]�X�5��<�FW3�\���b��R���(�����a��ضetȜ|��~��);��M�UqY�n��h⤺�V���U������51'f��<��<�L0�y� �p�U��Ϡ˿d���
�6%kά��2_��Zǀl���&��Ys����o��0�๲��j�PH�Ѵ�[��ģ6FS\�#fl��W��RʪniΊ�G+�LH.a�K0	����Xr
�
��|Q��U	���[�8�K���j����(4֩o-'�!rx�sl_uQ)�������T)�������Q�9$�P�Q�2�1�Iy)r%�7���LK�V�9�G, @鿪�x���^_�J�p�M�+�zy�8��������W_S�!�s�����hު��ݴ8hW3�Z_M��oRm`��Ι���f�\�Y%�[�{�L^Q�=WS{�lM<�V�i��2-;�z5�lW�5d���.^�@`�Q���(N���LE�!�_���DK_@�DJ 3:K(i�p�閔"�w���h�N��¥��u� ܉Lk5y&�@�"��UE2�l��;�J�c�߮�����t���V;�F���?�ں�yc`|bs�P��X'|aZ�T괒@�X$�s����v�����D��G�J�A� =���E���C�[�����&�@?Q^uhCJ}�����39�r$H�zF:��v	��*��z3y���F���A�)N �(�/�l���L�m'��֖z�h�i��6�(IX΋�����B{G�3>J!�.���p�d�����Ov�b��}��BHS�f�
z���#d��GjvZie�P��G�$E+<��r���Ia��hjYJ��h@S $|�m)MG�jay0l]ɻ�vdu$y�x�YI	{]��tY�f��a��)y8��2�խ&�OE%���~���:ͧpSs�c�������o'�6g�E�n���oI��}W�*��|�w�J��<35,N�M���O��J�%p�<T�����\c}T��(B�D�NѰ����t`��mػ}vmۆAj�}��dikM8~�8��&NF*c~!����&pqxS�s�d�غn��@4��F�kZ�� �|�������(�&6,�z������[ޡd\U��Ym{}��6�/���ڑ�Wߧ�H,�+��B�ߘ�q�Nl�.�nS7�<w��Q{��n� �5WȢN /�r���Q�Bl���v�q:Y�-d*Or����Y<W>���$�� ��h�<�N0i� S����"�{fM�wZ�6)nN��@,�h��\NYZ�T@"ּ%�M1��K�|�f�w�R�U��w����0\Hc)�@-5�4�Zr�EU��p_Y�W�N����T�3�i�m�Ҹf����*|Z��#��[ӑ���TUV�*�]����	��SV,-9�\^g�j�u�ْ`J �B<R'�F4NC!"/Z�5�ϲ>���:�7�z�G�B���z��yS��٪%^�Q�����=_(�D�\���g>X�Z�|`��x[�5�)�M��mEVV1���+�h��D9*բpug��L��ҩRɤM����4Q�@�~�T#��ػ4��	���!*U��Q�<-+�O݆�����iy�ɓuM�`=i^�����g�S#�z��bT���h�aݲM�W%��.5��~��?��Q��=zn��F.S��D�����TQ{����Y5�.[�R	i&��ض
\�����As8���$3�G0�o�5�JW����UيR^|`
���w����
��F���S��pE"!F�k��O� �c��ɦ+@Ok������8Fοj��I>=>�R6��d�TXDG36�p�u�}C6��⭷���n���b�4:�QW1Ҹ�DKoa�W��-7o��7���6tG)}��&����dJ�u0M4$d`cK��KN������QI�i�,m��S�K3�	,߸	,C<u�p�3��S�6i\$�>$2$`�O8�k��j����]y�s�s�{�"-!#�^bC$�)L�d�%2���05zr��q(f
��"'���8p�.���;�w�ND#A��Xq��5ѼF�^�O`!��Y_c]�Q,K������"��s#�]8?b�.����Uعc-Z�4 K���cע���s�V|���%9�z*��Ab	s���p]��r�.o:����~ܥ��v�3���ϓ,�a@JVP N%(��`��ɨ�,��O���%�P��d5�!��ڞ&�ۜ �	 �Z�^����z��s��r	ޛDs5\�2���s��˅Z�Ď�C�����p���̗�;`(�X$�P�K��dn
wT��Y~'G-uј�^L�8;���	T�'Q[�A=AK6�`ɥ}� F l$771A���]g�^�MSnvٹK��]F~��s����"�X�Zd�֡I+��W�[Y7�1�3�ʧ��-�%����x�B�'�3Oᤱ�"�L��e��<�7d�f��9x����H�:�	(�3�(�:!�h��� �OԀ�<���F.�"G�r6U��W<&	L�!�ŕJ��S�a��2Z{N�­DTQ7y�R&��L��+�r����'��!O�)C�k� 7l^�����r�,e���R��﫩^�P�
��i��bٴ�+1����;�˭RTLJX��0iZGNA)T�46Uc�֊�[Z$���b�u�G�]!��)mmq*b��[���\A<TG��
S̷���r��H�MwsLy*{y�5EM�P����d�m�r֥T�'xN]��%y[&����l7�I57ϼd�6|��Y&Ҵ�Dhj�d��?nM�!Za-T�z�n�ki�V��\���(f�e���:	_u���a����Ca�^A��6_k��8�o��9�����M�m®]���9���s�i��
Rg�0v��4(���@��dՇ�ؤ~+�>���x@S%N���sO�!���23���kFĠ��>#�D���T�LS�b�:��$�Ɯ�Hp��;�>jpZ �L ͓`��~c����!s1���4��}��_��m�p2f������h��K�j�>L�R�?e�}nr��=s
�����4
Db��*B��#m��G�W���>Z��Ăز~560�vwPӔJ]�ԞF
��+b�s/��?���)��X/2D�P��ܔ~��Y�Zg�2��5�ѱQl޲	�=�6�S
d\/��*х�2tZ��X߅L
�ݽ�w� C�O�Ⱥ�;	7����@~ճ��e���jckuv�?+�*3Q��gtx��$+��`�a�3���d{F-"硥R������ ��\x�����r)dR�r�(���-|5M�)���-B��J����s����G_W���S k���uT\Ԑ�	+�s1e�*г�S<(\�ڷ�i��/�m�טo%c���V����^��ZUPp��LS|U�5�^t��BO��6���N��1����r
��ۢ��TyL �
EA�\S2cR���hP���*�.i�����#��*��)i�N�@��뺏��o�`W������?R8�	r�GK<le��A>P]+�^�(��:Z��hr�,�U�Ȫ-�(L�l
G*����~K��@���^���,"��R�$}�Id��\ć�n���$铹�ץ@L�%sDk�*唣,Se�:rI��&�� w���w�s�[ �z>����
9v��y$	���8x��b�	ɐ��<y�,e�<��(ǖ�;���K��cj���5Y���Z$Um��qv���HoiZɤ�f��юpZ���<���0~
E�k��:%���2�S7��Q�����E3�lZ�������1���q*A�(,��z¾����Zn�J=��ً<&f	�5Dn�l�	���($/D&MQl"IAZW��˔U}��Ľ�C[��vZw1�^�MK����S&��B_wC+۱auvn��ֵ�����oB̓���'��:G0+!�������E*#rғ���2�I���-ڔ�^�E3-��Kgh����A�&��_"G�b�2���$D%����o�5�[������U��Y�0CڎHK&&'L�Id�P"���Ӱ��Bg�*/��T:;�-ڵ�OĤe�bҐx
������O�[���`�W�	�	a��!l��^����J��ui��l������a%��B-W�E6z�Ed��R�,CkLy	pZٸ�K ����׍��8�@]>��4���3^��Y���q������i�/\ı����W^�%����'�es�
��/1k:��u�v8�Q���
VWK�@�׊yd5{�˰��X�r��<7i�SS�8A�mC��C޷�$���~�Vx�����Xa�p�1O��KX`c:e��C�m֞��8��_K�h%�@SWF�Y�<��F�)~=TH��[�䏙#��:jUu�5����q�_>�*�D��E�խy|��fW+��G��%�W��ec�hqh�v��A�	$f&4���z9�S�*�K�W����DR�3�Ӕ�=1�F�T0��-Ъ�vO-�^β�3L4��i�*t�B͉�4��#O���Η��R�۱%;����'�Zh1ң Q!��=�sU
Y���z��HZ!�C%Ӽ�h�Y�6�I	���1��s��YS���}�
�ǆQ#���R�m�����E_�b�2-Z�;�)���["������03s���
BK�;�'�&�|�z۽رy =m!
Y�f)C����ر��RE�n~nκ�^e9��V�l"$ʳ�7��΋����,79��ڜ�_E��b��d����r������ށC� ��Ķ�^�����@2O�h�n��?(���\b���VeIkK�r����M�!F��#��S�EI��+߈
�%������?�u+cX��Jҙ�8����+�m�b��k��u`�� ��0;~��*��ҏ��;q˾�X�Ků-h�V�S�������8�c�߱C��ӧ���i��"e�J�}��x�\�{6���m��r�q�la>�B.Z�tD��
VѼC*-�tɺ���2FRL@g�xт�u)���'�e=��~N<���0�Yf�)��y�}�E�?~����ϟ6����:���Q���芅�dIG�G�vS��05Iz$��U�=�mx���R��������ixÝ��Z11>eD)1#᥹v���\�$�\ΉB���O���fL��=Yv���[(�S��-�0�ұ��D��dM^<	W���<��Xx'�n�y,L5�I����*N�b���h�DO��A��@��o�0r�ZM-�M��`���

f�0K��BW!r�@E��4CCk�g�uvQ,��^>�2�_:���6j�*�p�z���r�Q����Xv���P~�8y
	j-��k�$Y_)�[^uD�J-� �����(��PА�z��18�,�܌5��JEڦc	;��9�|�AV�~�*��ʳ6����]%=�B����;.�伿��*Z˲�=	b�RƸ9��7��=Z�:<˓ś�(��q(�JN	��=��a��1ֽ�8����Yj�]����q��Y2�"�R�}����@)�����Z����5xh�/-�S
�[��J`�RTD�0��ݻ��#瑘��G��0w�L:�P~*?�Yh��mX�ʯ�~	Z%�H�;KA,��F����P�{�<��,2�G|g��ؗ��5�&�O!/����"}�X�*�	R����p�����#�Sk�,�_���85{�W`�(���4��$m�ϖ�(.�;e֫z�"a�Gݏ�^�lX���1,L������Z�i�"�J���rز�+{[�d���#���SϢ��QުU���33��0L�l3S�.Yo���s������!��[��陙+ݚ�+��>s�_y���@������	���Gڱ>F��s#I�Q$�^m6Q	�
cf�uSj�Oq!�.�ފ��X��N�l���ZV	�S�}�j�v��y��u��r`n>�wܰ�ܸwچ�9�[qp�z�嶍���M���܎�ن�;�c�����v��q۵�q��m8�vn"��Z����Z��]���u�m�:~k3n�an�a'�߿������]7l��]��o�*\C�����a�V��{���}�f�zx�^���h�, 7Mkx��u���E�c���J�P����a$)'�y,�]���E��	��%����%��<��R�41	��]8@�%Ϫ��դ�|�$�1z���&��Ip��&�f?n��:�ZM���l���IZ�Ā��ƺ[�Yx����{�H����3G���+�E���c��8 E	���P�hbSTi�ߐ̮�Zij�o'�O�P�J�-�
q�jcԦ���*(�t˾��`�'P#���� oYk�WgkX�����2�-[�hy��6�h���^�+dtfA2A�X��Bq���g)H���� -@o�SB�&{��V�@_W�r�-�h�{g`^���5����l]���~��}�A6��α�(cJ�B�����?�4Eᠱ���nlڲ�3�tq�����xv�ڋb��F�O�����~_�d=�|�@kA��!�	`%f���0�ZA�Q#t�@��a��(/)����g�	��X��	�KL���y�G^�u�_`�r��L��L��9��v� I9�߬��!w�6�������Eq)L*Oę8]d��'1OU����ق��S�ҥ��P/j(*c.�,A��F���L�<��G��獶�m5�$����<�o���:�ઇ_��bX�3���Vӳ�/N�G`��i$�'(���O��g�0wV�Z�S��{�@�Ç��M�mZ�9]ֲ:Ba�Oީr:@�&#Q���̺�.U�����p��7�r`c���8�j/ҋ�F)E��_>�`�f�Z�l��t��A9�X���%�ىD6��YZRy�i�YK~�py	��ZO���F)E%1�Dk'[B<Ҏ��6�\<Oe,i^��6�<#�0�>
����4n9��߽�\�V�<�]x��g�ģO������T�y
��}sӴX��3r<������J%.��_G*�6�SPf���+S��r�?��{�)��������Lg#_�:�,E�a-2�GN����{�P��n�i�+0E;���Ĉ�EW.�~�x�X�<��M^tv���1�����_x?~���Mۻ��?��AZK>����^�4cEw �7vb�@Ȣ�����(��7{Z�غ�C=q��<��fkw�k�C"��Ԇ���ysh�u�Y���!�;�-k��.�0j��V������xOKk���E|�o��z�_ug�%�i�*Z�EZh3��TJF;�^2������PY򠯧���j�*(a��Sa�D�mT@h����� j�/3�Q�2��P�D�!yϼ�����}X=���`݊��<�;3�D��z_���nؿ�y�7����%��҉Q?7E��$qi��q2��@�B�G���1�=�(���JUw�i,��(�>���"�5۸V�T� �G�Wb�2����w�Ӻ4���3��o菂H����[̬��Ž����Jd�TY�9�^2Ӓ�R7fR�E����A~��o��i̞ݡ2>�� ��ZA�fx��r��F�)��Z�N���E$�f�(l����%!䣕0L�Q�3u�9r/~ei�ltu����w7����D�a���%
�&r��l���BЃ��X�f5�
�(Ҵ��Ӽ�m ��ظF]�l� _G+�Ԏ�?�ԨC�YmW,<։���ܢ;JZ�@ !�|�X���bӤq�+�?�Zj��EI9���N{�y��h(R�պ�'ڽ��J�/<s
��gR7�PK�i�J`4S�ŭ	�r,�PQ�`���P㚴|��E+��c�4�<�AJBPc����0u�&�j��i2��E���B$�H�t�q�%�-S�S�Ԙ�����̤u����*��TtJJPѩ�I�ZuD��Թ׊ ��+KK��41�
5��_&O�rU��J����4]E�Pσsg�j�.)"nYJ|��o��zbu�e��@�Yޘ�����D�ZC\S��Ūg��ɒ~r�')�f!��9w�\lG�f~n�2y��I�������L�L9�h}i�%��-S��N�b��>Z++d�������cx���(���z����g3��F0�b�[[�Cppp�-K����,��
�tcRvI��y��C!D#�
_f��������݋��8}�.\����~��z�(�E������<��8��-(�*��z[��U����v�X'r%���B����Z��N�;x���\+S��)3�'M�Q�4�)�ڳ.ͯ���`�0������d����y���~7�z�צWT���}��л�����l�4�?�����G_@&5O�g=mѰ�i�<�|�Y�>�z��!�Wsp�{�D���#ȌhW�G�d,i�%A��d�N�w�%W~4f��性h[����S�N����̻�V�H,�q���lN��@�&Z���9�h~N���˧�m�����665�<ɽ]:vт�6/Qx��$�VQ�5~P���/WU��ֵ��4*�l�r!M���!���BFu�U�7Ѕ�X��dD���VV���s���tK��@Zz��2Y��ژ�"K�����f��0�S}�Ix�ؽ��6�2�S̳�VZ�*"!���q�����$f�P�e�Uf���9,.�l�5�ˣ������N����?�d&I�K�]�*?�Ra��W!�9��'-�F�A���5o%mVcw� ���1���9����q�����'�5O�j[�
��>*�uY�R TV!L�W�.MP�����%��'"Ԃ�
�%8��HJ�ە�"���)U�Q�f�ڋ�gZ���Ҹt�͆`��JŞ�m�m�≇_E���:J��:�r"��_���
r�$��dʂ��L����Yj�2�V�H����ͫ��{	3����PcҘ�:�ޥ��L�W�r�$�<*-��i%1c,&�h��:|�_br@������A��O��Ͻ���.��"�H=&�
Y��L�C�B���8��m��(|���8k����e@fm�
��]�j_��ښ�+��%p��H�"Y�
Z��7�͸D-?�u�ʚ "|�妉�n*�l-D,0W]˙Kʟ�
�5�\����%)Uv�]�"�R"�M|�rT�iU��X���
��1�Ϗ���^�Z�v�܆�n���#����ס��ێ5�AC)�-mT�[�M�T(u��aE��{i����8�?`=*/��n3�r۶ho�«ǎ����^�ݳm-���<M�x��H�9���G��u��*�h.�͏Ӑi�H���HUc.�"��Υ,^��)ohH�P��^��1:]¥�,*��D~	��&�K���X
�g
�X(#Yt!C�K����<Fg�+`>]A�@�*�"�g�E�Neq~t��Na!K����9���.���)*,g2S�eL>/Q�[���O���6��:Sx/МH���O,����P�K��6g%����<[�f�[�L����;�b�U����؎��W����7�nj�u�'��CAlپ	�t	/���D�tM��������HWZ�@�O�ܶ<�ّs�^�O�1�Z��@� ��̃'��C�q�m���C�q��شf kV�b5M�4���و��֓��9C�,���4�>4�F+fE�uiJ�9���bܫ+��P��[���kZk/C-E�i�yi�nbVsT�u��֙������3�_��n/n_��hӣ���� ��]j�$G�X$@M0�k�v)��U(� ��Ծ}�(�صg/zzzqa�2G��LG��V���'��� �2�A���Kd1�^���;H*d���L,.�908�H�3󘙣J�*j�]V�r]�+G�[�X��֢��2E]#��TsΤe�ةKS��Ѫ}��<?5��s[؋(��OXK�f�6S��#�$r�l�� T�p���H�<a������Fo�P�1�x�$�8�KJ���ŤU�%�mqa2��C����u��b=8`�	�R����4�QV��V1��Xb+A���(����T��mˬP�t,��'��U�=5�M��ջ՝�15}��.�0k(\��(��R�� �����/VZ�P����3&5��MeSn����?���^\��s�u��;��q���#ۗ����`Qw/�&�P bU��w�a1o�.�k�DYn�����ҥ����ƪ�H�
��s�z�`��ؽn�����5��J���OԆ�V����E)�r]ה�1t��s� :bDv���n��{�H�±�{�[�o���b��^�	=��d5�ò�uv�� ��.byM�#:��=�@�xA����P4-�G�2����S8q���"vd�Y.J��D�J�"f�TD�=(P� *��!�JhSS�z�]��޲d��bl*⎛�aͪV�1����4�����{�~�$�Z�cϏ���������E|�����_���x���c��0����3�������{�}�4����rn
>y�~�(��ݧ���?��>qO�x����_�CO�·:���3��<�����y=qO<����ֶ����S�q�ŗl*���
��ҩ��IM$��X4~�)��@�3��vf�<w�Y����[��u%�e:Mc�EXe�)	H��Z��H�����n[h��޻�t��1�P$x��o�nx���PW�V��u�Tv���;���q�N�dIm9d.a��>|�}����X;Ԋ5C�غi%��ހk�ن���x-vR[S,�ŹIc���,����||�
<�?�CM���4���M�p��<��F��q�..y���ҬMP#�����ji�6�ϳ���0�ʓ(O��m��b;���1�/����F_o��M��[���Y�DK�
"�B���
�oi'qt���X9���.\<O�m>��d@O0�&mr�����5c-��>�j��{��q;��;6+6`k��R��	�753�9Z�D��V��!KC̯-/B"�u�[72��RW��Z#9�Z]�'[YV�ui�R�L(�� ���@�S>�
.~�_=�Q�ir��Ŵs�Լ�$r��^�@����̼vΪKSV"��W$�?��1[��L���µn��F����na�H[�����F��t�Pn"�,r��%��M�&XӺ��FM�َʋ��݋.�y���� Z�Ukũ�49]Qs$��]�ZZ�8P㘬0�3٘4�(oJY*���c�r��х��L��v�Sy��}���侽۰je/:I6��6b�`�1�og�l/#�"��b>��uu3�2;(T�/���q�R?� R�z*��O�,��zTY6���TgԶ�K�)),�����}4�?D5�V����V�	.,����nZ8Ŵ�uG�1���������ɿk�j����K�m�H�P]�sϝ������a求.��k!R>�/����%�V�L���#KD�s���ҩJ�9a�h�MMR��y-��H�g�^0k��o�oJ����W��ዘH�M�o/�/�E�W�y�^���ֻI3D�s�R�z�@��q-�H�|o��0B+�;�D%d���L#��.�1��a���Had�$�>L%�py6���Kʹ��H�HU�X��q��(.M$19_D��s�V�`&U����Ӹ0��UX$�7[x1�V15����˸pr۽c�BN�8�W^>²�_Ǚ��XG-��E�R݊n���u�+�=*��A�E9	�4�z5��X]���"~%l��~���}Tx�NE��I+�궝;P�^���0����m��x�5�1�J����}��rf��8?��Ӈ�"�N-'�br��fP�M�Z@��ş�u�6����V�%�H�ҏsɬ-I ���&���믥e���gP�����տ�b�л���7��e*�Q)A�Z�Y1������,zV��j�dJ��-��^�DT�L30�[B���I��09��/?��hw\�ޥ9������%p���m[�H��՗_�5�r
�Z�R�Y�7݈(��\u#�,`z>�i������"F�Fq��)L.��(�����Z��y�!��(LU@���[06N��s����s��U���Ƣ��@�x�.�O�=���~��4��<��,"���&�u��=}�[3�4�A���<k%�7�~��
�I�H�-�C_�	ï���G���HM]Bz����O�cjd�m}پ���H,B��9�X�Q	7a��Tե�6���^^W�Vj)%~�%��c�����1��J���a
h�0��ww���=�ű�m%H��-]�B�m�-X�׍��6]�H+�F��n=�e`~D�>	y-�[]�cV����b5� 
]��
���DPQף4�*��4�V)���lc)S&�K(�=Z��˖ػm����[bώx��w�C�w�q��|-�� n�y�ٻ{wnƎ��}�*l۴�vo��7��-L7څ���kv�[o�=w܊;)�wl�D~�a���y{�R�!-T�,�Y��g����ivU�>�R��Ń������}��-h�Z�\�	.� �%����<N� �炱��΄���nd���$�{�HS�i<Xc��[	=ma\O��
R���QG^>�'�|��,����[��p���9s�)���5nw��	{�U��
!`J�:y�<6���1Z�Y�^����\��W_}+WR�����=fNO�H��{�9I�R �o=v_��s�z�(�����+�c��x�ڦ����ս������-��,
�)�<U��]���5�P�ͯ|�	�*4@���6�PuG���uXGc�*[ĳ�gj�E�UC|Q�y��/�Wq;�1�{���\z��{�ǲz=E���B�W����ͤ��t	�7���ۄ��)���h�R O��9��]`]�)����H��5�P����lVJjCYi�Y�ڳU�%���"��	Ǔ�f�z'�w�,���F.N��
X�c��>=�����x�w^�q��=��
��5^��#�4ֈG���sǍذ�>W�c3���|�����?I��y<��sx��q��(��݇p��bC���m�����OZ)�>V,�2�b���`�i{N��zs�9����e&S�3�n���:�~rGkp~s���i=��P/,!�(�؜-�H�E��
�����F0�m��2���HgQ,���u�Vt�*u�ԅ��)�]�Z-�r	2k��� �ӊU�6�s�*��+0E
�,���_Kw'�m-��
Vj1TpX�̳��ڶ�R+�0�x��ذn�x'Q�CX�'�D�3p/�Q�9UJa�k��U��q���0"<f���ұW����E�W޶L��j��r�Q
�Kǎ��H�5��0ԶW�e#���D1�$dR8&&T��u�ytqMp$)b���\#��^��U��r{,nˏh�s�Iːhb���h�S'�s��A�a������LA�	�5�ߣ��T�Z�$�E#�����f�SR�nM����uY$�T̓��Ų*�uAև���e?~��ǟ��o��?�>�܍�㖝��F���ƪ�v�S@vS�GٶZqDz��O�1�^�u���V	x���
�Ķ�+�c�vo>�?��7�/����?z ������v`Uw��]��"�W�ֳ6��^Ji�5V�M�Na�eL�nf���g�*B�O���*�I��9�R�7
ty��ca'^��sT=�hzZؽ��J0y@Ǝ��2�C�@৩hu�Q'�ɒ�1;;O0Jb�<��#ѵ���|:)Q����#��7���|���������/|���G}����_��_�o��o��'��׾�^x?�0�������_�_�ş�_�"���+�;a�)	h�S
s����^[,�bևXJs�W�r�'�a�����Ci�"�DH�.ޣ9��Jq�<�_���}ze�x}~�JW��AHK_i}Ś�<o�=rvssO0�բ1R�k�r�`L
V�,s�E��<'۾��9��A� ���|��f+0(/u����]�������-o{�7@c��W�͗T������ ��Q��KI�e�{T�-J]�>���m�M�����ƕE�g�½#�e�#��Q��m��[NI�?�E�W�<�xE-U�໩�<�X���)�^ޥ¸*�\ٸ��lۼ���u��.�����.����G|��<�^:z��{�_��Hp���'�郔�l|Ͼ�;YC|�"����!}l���m̜̲7l*`c����l

p���*Eω�$|ihi�B��L2IY��g��L%�\%��XA+�ì�T��t1�L�E�X5����N�YM��B���D��w���w�*t�ZV�@x��U��v�sh*R�Rd�:W�����o�5��E6�����ĺ���Ƽ��8v�$5�ftuu����T)�^K<n��n�4#�U �8��%y|���n�W���CO��D`�vO����/b��S����u)��ZY���B��D��I�}�y�^�����D�C�N;\��M��&�^���@���GlLPq"�,D������&~7�xKT7Cc7��4��PPk^�C]]U���w���YVK��b@V��bj��I�E�,%���(���Y�
��n)���4�V��!C�E��z[q�M��O�������g?���~�~�l۲
!
D�qy�U�fS��@�L��z�Gl<M�r^K�8�<:YW�2���^%M.�l���Z�ؿsA�;���[���O������b��6�EU���F`=|��Fa����7�l�a�YG���HDRr*T�*��i�(j��K��4V��	:�zY�R2)�i�)� .F�.��І��gӀ��*�wu�J!�XlooZ)��9r��Ä�3�N�\�X�.Z��	2qVPb�ݽ��[���)pT���*`v�؁/|�wmi�*�XK�i����bt�ԅ�$�|VєB�
[���[,�g{R�#9h\N��q?�a*�b�����A%H��*|��m�`-�i7lC"�C4̪1#@��m �P+�2ɚ��(_��&Ґ��H�]p�ey�[l7%)��]�s���,�5�ܴ�X/e�]�=�J���Fk.L��|tI��-T�R
4��JV����;4$�uO�|��*�I�&�o�Y�
�v��!+]���)ݫ�1T�׫��f�_�ڑWM�H�G�e��eWY-O��y�р��fᚙ��Q����Rc��G/M���z�V��~'>���`��m8wn�S	�:{	�s)�J0�:s��Y�Y�iw��&�=~K�~��@1�1m��=��x�*�VqPƖ���Cx��VG0Ph��fqnn�khh-+�	�)�k�riڧJ5̧��SSj���f�ډ���������Po�E�M�N ���p��7c�7`p�&lހ���m����P�l�5c�~5���!�(�B-qh0������������W���<�۟�5�P�fY兙f�"ΘБ+� @nm����B��7��e�9����Ԧ��9;��[�i^�����VG�0N��C�bK��i�k�)ds�CZ;
N	���$fΞAjj����!����Wor[V�.��'�n�"�o�,�(�
�8��%���%Z�,��T�S�G��FU��Ҫ�1�P��d6�U(h*&`93O�����wI�/)���cZ��	��GB�v�d��+{q�{񱏼_�O�������/����޷݉��Z<�&~g~j��{֨8���M�s�%
�J��E�K�]���4���U&�RToω���R���C��|?��,�r>E��#����:�א�Њ(>���?��������߅u�[���;�@0�Z��`�Or���pS�gu����Yg
��R�����z�OW�%fff�f��I�Au7���1����R��Xi�:�Nc�G{Ѱ�U�?����ԍ�$��&��[�~�)�|�e��Vb;�;
��~�f<t�"]�x���O}�Cx���a�e�N�0Eh����{q�J�h�rG��<H����u�˱B4kʎP��D�8�B�ۍ��φ t�HR��<�y�e�8]�aJsEE�
W8K�<q�,R�*�����HTc���b�ߑ�'(�9w-G�̰�iA.Qa���s噸o�U]IX4�����r_O3�H?�g�Y[L�L(�&��yNQ_<5ͩ���-/i�� ��X0L+�FK2�l2Mj�a(u[Z`��,���.���Z�4�"����bpŠy��t����]�L]]���z����
2._Yh��+\֯��jl�wS�ɑ/���hxo.��P*�M����Z���۟����.5���9<t�·!	���)ؚQ��mk1�ׅ��^x�0^z�UZ7at�u�曯Ê�v�9;�^83�:�����jM?�	�����@�D�e}�A$2r
����6�$���<��&fX�J:��Ʀc-�n���>����6O╕��z�  ��IDAT\��QBw�,�&,�XGS����S�`��t��]̂�H�OQ�WP�,l��@����ȩ�}+�i�.9u�'fؠ�p�Z7�a%Z�{���,S�{؀
�� @�V� g���i��j�=�+0C�ajz�DG�& ��2�����9{��$���Hg�5���,-�Q�_	9Z��6�l��萅JQH&r�H��tbݶ�Hj�+2��B��`�c�ّ��RG(H!C��O�1u���R(��Y&Z35j����R�Z�a2,�T�C�#����X"��V`�[�NK�Q�Lh��d�C!����ŧOc!G�DY��l�$`I2��o��>M��I���N�C�:Z\��-Z)��Kfh�EJ��YK%Y,ܔܴ���n
/i����A��-ggY�sص{����?q;�?�k���E֨�
�sl�E�4ՠ&m�����X	�F�v�y�|�IĈ�뤺�X"�H;V�Hn��|��zN�-Oa����X\�+�$�S���®훱��=�u(:�t� �b^�O��~Ӟu�L�"k8��#պ)�Kl�Z�`A� OQ�f/���ꊧ�('_�f(��;i��VF�ز�<#oYM�76�gWK���HJ"�P)���N�����l߾� D+�K@jQ�0�%�./yPk���-[��} �^s-˻[�n�e�ԣp��1����k����n�l�FSN�
�|��]F�86��/����R��Aˋ�	�,��y�����Z��E�lf�@�;�4֬��M��|O�ό��gaɋ&ZU�(�@�5���֔�U���L������L1]e���vn�Bi��jOZ�j'��
�ǰ��z����	x>���4LvnY������.�9�����Eh<�|��(��iE��	����KF���s�.|�#?����n�	��r�z��m�r���{�q+��6,l�.�Yݰ=�[�����O�؁Y��L��HQyq���h��dB;Ҏ��4h�,(*��5=y��KK�HR#Y�I�1��-�� i�BN�����������E�ܹ���O����Җ�i�PS�!�R�
S�L�h3����:������~j����&�;hܹ|��$!f���A���>2K�@�� ޳�b*��ѳ	?7�LA"E�ֱ�R0�
fg�0|��ԥ����Z;�xh��`6I�&a�I@E����5H�D�(H�ݸni����ҙ3�����իѺz%\�d�N���E����WP0�169������{'��L`�D&�6G��jY��9]KT��[J�*Ҡ͚R}05�ة�FM�<�۽s�:͕��ɺ��*]��OxzI�A��qY*e�:��qbl��X�)(�Ӧ��F���kZ]����V��(cX��6>�`s��vԣ=�{�Q�Q�uB�%29LS�ұ;����j�|O�<%���"i'@���慩�E��5��\&�tT�s�r��i����D$ɑ>s�g��7�����9���N��icYIO�V)�%�I0i��@�eъ��j`�2��5�.�V�����ZDʈ�F�.#i�_H���&��v����AӘ�j��Ľ�n}|j��# ��h�m�����O���=x�]�aת64e�h�-�'iuj�r�oS����sQ �>�����.c)5J��D�����,��z�Z1^�4��+�1Ŷ(�4��K�\ThrK�
Tx<�fe�m]�Z�@!�<��T��v�l�2��S�W��<�=ZhY��Y�Dc>�.]�W���8y�i��<�}��>���/bfv����1���|�qq�u��-m���f���\^��޳�p�$�q`n���,y�61i~h2[��,��iC-ҍj��Y�0.�=��y�u2����C{�*�ύ��P�k�#hƚ^Z�uZh�qT����=GД���<�zaK��ɶ
Vg��\D=s��Σ�F5w��IvM�qx|.>�@n^�.�ݪ�'�L�9?_a��:7��./���3��b�$�i��
'oPa�<�2��Ŕ3�U�<c�5-zOɻ}��2�2I1m���#,w��Ɓ��q��7�'��&��o�6*�z�m *��'Z�k�v�1)�F�T���)G$M�jrk
e���<&S�"��ϗJ��?Q7�� V�FOC.
�r݇�T��B��~�t���_�(�����;bp���M����];��w��V_/��-mݨ��l�ԚXi�f��1ĜH#�"�<h��R����R[-3�ʼ�1���wZ���m��t��_��,S���h�v+aab���������x��:�@�&d+-H�$�.d���5�8jT]���Ԉ�eU��b�Z��SԘ�ɰ�S�YNa��B5��w���CKL��yL^:�J:�0�������Ato݈���(�ȩb�@G��h7-�`�r�K�N����'^��/`��+X���J�¨���� 'h��+
 k|V��ް�?�����Z�,
SY�5V��ޤ�ٴ(\$bկ�$l\Lj'}����кPC���a�BV�jCu�^��{r��������*T�H)T9�X�GP��,�H[�Z�#�5��}�hE�	tU
KMuQ�3��Ҽ��"3�z�A�КSpe�y�n�<�I*
�FE&��d$���*�_��-w݌��>���|����ᾛ6 �L�\�F�Elk���J�PPo�Bg�+K͊����2c>d�QhLI�j��y?�>�\�x����,�����-��csj�t�R�)�8�0��V��k��g.Z��̡� DCa>2�ރ;��{3~����ݫr���/�7��B�ڤ�I�w]�VE3�6��"D��ɌÝ��Ţa��4�g�ws��``�>\X�K2_>�#lZ:�6*��'���H�HJ���4�gfx=�
��UC�6�KS��3��u5K`��������A�l�֬]�7Z7���
�x���ho����"�iM�]�1��U�===oޙ�×-���ӱU	���-OQ뺉ʅl��b�df�,��߶��^Zi����#O�y.Y ���-�h4z�z��RI�A!�T H͡�� _r��$"�Ex	Du�R�4� 7%.#q�e�/���G��]��:Me��8���e*$�s%P?�Ĺ�P9���� }�	L��N<J%���)��"�s�"��cT�^�{͡vS���B���@,��Q!��>�^6��<o���R�����~E�r��X��{h=�f076���g�]�"u�ȟ����9��gYt��GZ�f5�Z%�J��^���Hݳ�Ѩ��&�(WHx~�{lL�[R  ��G��ICm!KZ�E����o�'��h�u�`Ǯ�x�{ދ�7�E���x:�ڰf�*�z��ذn�ቓS��) PDUN�e�g��v/3�~����Im����d�8�g_���7�tEc;�V�l�����\�4�c'���#�0ryssyVn�����6���#��!�LA7��V�zD�%�EF�h8?ț��O�`jwws�ܡ/�?���-C;�r���ش~���,�Q?-;iTY>K��:�s�z�߰���c��t�G��T�P�7��P�l��M� 3��<�ӫ71�ۤ@8�S)�� 5�r��"K'���$�ܭ�+��a�'��DZb�Vi��B�֟m��3o�&
�b�	�.&�LΣHeIn�Z���#h�Y.	Zu��:kbR��Ɨ��9�*�`��q�a�V4vP4G�pЃtz���b�L�w�]T7��!�������kI,Nc���3�{����[�|'6�_I t,R�z��ܮ>�jɋL]���h-m���E�`�MJ�~��Rxk�Ȭs��hWʚ�h�9Y�W�ȯ�=���גc��KT��#�]�O]�����M7݈��������+�iUW�T&�K����X��WU&��O��MNA5�$h)�&
Ds��Li"���S����'1�I�i%9)O�TX�,��M�R'�x�� ��hո��=�!Xj(D�t4�Ou�)lU����m��џ��qǝ�I��Сp��𖷼��v�t���'>�����&PUߪ	�*+����|�J��ض��o�k~�څyr/wǞ8��BN�O�I,����&�VM�'����W'�7���Qc��F��C�̺>%�5���/�����<��/յ��M)�Ƣ�z.�@���W�Cz����l� ���w�hy�PY�q�/_Bw<�{o?���]���~'>�3��������ޅ.�R��J~��C�`Z�֫�N�!� ��H�0�;Qtk^�%M}1b3�h$=[�}��OSN>ZtW���
�;����8sHa{�%�[㶊2%�]�zj+�E:/�ŧ����j�|�i��͒�w��j�#H^I�Y���H�/&�I-�^w#�����0��⦳y��S�(�AYfMt��e�ׄm[�l��ҥy<��8r�U:��5���-��,��(*<o�3a�dEP��MBB ��r�{��޷|����o*�I��6�W�ǼV$%'�|}B���i�j.J�Zs�Pg'5���$Ο��4�M�M&��\�`�RUģ^���8w�8Ν>n�Y	��Y�H��]A�V�hĲu���S'q��I�t	�}�馦H��0�BS3mc��& ������F_3�G[ԇ�@wV��@WP����*�Y�1�|�&P)�To�e�yb=i�#��u��:A��V~i�y���~5I k/�b"53�����2[��Т%uT��5V�աe6��±�Q�,V�t�%�Aqa��1TSh.��_ʣNЊy��E���Fjv����M�,��(�
���7Ri(SP����:ͧ�����&�k.��65��5��Zq�m���(~��&(��$�Tr���b��1#�#��@IL/0R_�4d 攃�6ugj�Ht�v-�ML��kVO�S)��"�N�~ޯ��:�ѱ�/��d|Kg�+�jQ����M�NmkC$�"�*��P���g;oٲ�����O�o{����!�c�������:�u��rE'�?�V�0�-�D]��O��zR���4�ny&��Ifҕ����E��c-8|�2�|a� ��I�_C*�r�Ch�^I����+�X�hV��h���p4n�[Ǐÿ��?��������������~�������sZ1�L~l�(�G�4�r���w��� �0���#O��s��i_�޳H�	���B�V�=
�L�|A0 ��'��՚x(*������Z�D�����zr��P�W;MOMC+H�j�_�
��8�!;?���E\�m����~����ޏ�;��n	��� yP�V�s�x��w�_����O _�O?����O����I|�ww�r���P^��k�a�7Pq%�9�2-�K`{V�m�W)^*ѣV}׾������i\����"�#ڄ��|��+�B�Py�qrы<W��f���ynJ��Y��&����f��9�T��id��_��<Aş2EX�VD����P�MͲ�0���G. �B8����o�{6��@��Y62�95�Gy3�� ����r�z�	�z�(Z�z��������y�0�N�&�����lU�Tj=��X�q�eHs/`bU.�l�^ڮ:��<
��bn�4��Q�K��z���$�3�|��V�si��i�/�G��֘����L���݈�h�ın�lX��P9����g�[���(<i��hRO�MZt�Z�L��1�?w�VX���e]6Y�Yu�i!X5☜P	fm-q�]��9[���X؍]�Vb�@+.���9�gYnj�6����@��S;�w�a�G5E�M�RPh���r�����!��ͩ[��GAD@Qčz��x�D�˚��uK��\4uQ�S�5�ȱvL�h&-4y�����H󛚮-�n߲1 �����Jغ1���\8%'�6�[Gf�a�mcn��f�B[��i��Z�ݭZ��4����n���TP(\eՆ������<�3A-�q�w3�r�V�p�8�T�#�������x�O�����Gc{�ddMRp�~Ѩ�|M�q�U�U��69�H;���PI*cd��Ɍ��p D� B���ڌ(@̲�M�n��TMY�+��p�i�%Yʫ~%�~	�!�l�<c7n�7����6�LexMmǗ�9��V�0+�Y���䣱
k�C�� �o�v�S>d�t��LS>�����,��K��Znv����r0.|�߷�4Z>
��+�z�z�^>o�����Y�E<4�
C�V������V\{�Z�ر�n��]w=�nق�+�裏���W�E� @Pa�DZ�vbn!��k7��<ȗjx��9��<>��GN�+�y��)+�[����Ku�NKJ���(pl� \g[6Q�h��K��m_��.`��.�ܲ�V�ƹj8|��7�`�%Z�
è���Ĭ)��x�-x���ƶk�e�5ɚ�^x�Y�$T�j
׮�o��'q�]�ؖ~ʨ�9�iI�L��ap�ߔN-�T��)�C*3�b.E�Չ7�}��Y�:y�u1�(����6S���>��m��&�{���K{v�����|�t��X=���C�R��W��9*�6&����~�~���:5����ܨW��k�a�4Z�x��(.MQA�2�����!��'�HLm)���sEd��[�@��`�v?5?������S��	<��s�򗿌��˿�L��η�����O?cs��f�J� ��$#'#�j
4��b���0�?'?��?�Q�9���{�l|!�ɫH_�Zy��S�`�_�!�l�v$i�-Ȉ��d�e�6��Cr>CF�cߞk����g>�}��ق�#��G^�1��=ضqn�~?6oX�)��K#�O٤˾�^(����85��Y����Ep,�����=u�R�Sx�j���jf�Ƒ���r$>-c$OD�F�e�V��(��� �� ; G^-W���ol&�yPW�R����.��uD� ���s-[y��lZ�L"��֝�p�w���"M!j��?b��JPa�vZ��ȓ҂+���7�S��@�Da������ڂ�.Zݚo�{��Y���EG)�IW,�/i�
�	��.MZ�9��*ɓ�٫�M�>���Ǟ]�(����5��*�7��G���ջpe�q���iP�b�.Z�g��ad��rS+9���Ճ!��$YN���5�/�j��T��	�v%�K��`^���|N����Uq������V���
d+y�Q1�u�3g7囿��'+�]�{|���~IXBWw;�VX�au1ի���)	���#��܁nT\��h��?��h���`�<��!����jh�M`M�r�@�e�{�����>��/�_��W�ϴ�z�)|�;�����-��g|�_��O=�o�~��Q	UO������!��H��(J-m�(�B�����#O�B�ڋP��`*��l*k�׮Y����q���c}*nf�U�bg=�/�iL�@��oNM��m�U�j#PW�h%)>�T��M�W ����o������ƃ;Q�U������%�Ơ�UyZzZ�����ܴ� �9�ZM=Z)^�ʻ���~}>��w�k�0lO��M�g
�{�>l��k#�P��L�y5�7���U���Cc�~�����<H�$�w4X,�"&�JaS{�����f)����hZ�d=)�T�<d��X����;$܈�^&0�ܻ?��O?� �%Zxr�|��s$�D����Ȍ��
���{'~��߃��?��[vP{����7m܄�CC����Y�oơC��[o�M�ގ�;wcϵ�3�!�:}f�B_����$
d���sڶ�&cj]5U�ZR�n4���a���*�ڧ^�,��JW���gN]�B5�{U��gdq���!	k6i���蘍=I�X^c��d,��䪺!!)x�x����盚�V�޽{n��-}t��0e� �N�{��^z�9�?oV�����vӎ4���'5������I3ˢ���ML��S��Km��KcǦ!|��ņë��J��������UVQ�5�RS'���;vy���p� Q�Š���X�Ҭ���_�i��ml�����b�j��V��c��-&��p	M�A
-j�|�B�g�>^w(Uˬ;��3��l�'}�]o&�ɕ�LM��mPǩ㗭;Bn��yL��%5p�����e�#l��Ǐ��+��2�HSn�M�m4U�0u�ܩ��a���eS�("J շ+D�G�=����5�A��(+ꎑggP���L`�I���G����b��e�����(�Ȥf��É,$�\�LuY:VYc�;uɺ�x�d5�ل_nQ�Kc�2{��R;�U}e܃ɱ�$!�g�N���x����~�W+���[n0W)t�t�B��,-,Z�3�,6���)���مEZ0�ho��WKHS�s7��	ű�	S�����RM+�4��{o��ݸ|�"J�QMX�����x���Y�
R�E�Ck�Q�`�$n$?�ٽ���Y�9����h���B+l��왳�Fc�5'��s��������0����f^�'���(@��_��-*�H��s*yny S;sS�R����_f٫6n�D�E<d�z(r�Y�L��ߝC);��Vn��:*�����cT��N�)ԃL%��;_(���Q��>�_��O��#���(８�T�O_{���m㉱H���򱏾z�=�%�e�Py��r~��KNs�x�T��H-������,�/]F$ގ�t"��<u����J^�㯼�s���L9�����FP��j�C��f�vRA�j=�
�N]���T�g����&�����y�9�2������3���?u����1OR�¤�W�����T���#�4�Ez���U�+GF�l~�����m�N��o2®ݛ��3��p,��h���"X���Ww�8�m�E��6~�5�����[Ȩ
hՆ�jPSߑ�n5�H��k��i�7-k*oܤ[������Ȱ�5�Ć/��m �{M�At
VݯN0학J�H�"����g���*��[񎷽�����Ncqf	Z��Bj���"\�8X��V��I�eR�uW �)��,<��=MP-�	~�*���&�L�4����Ed�B��V��p��E���A��n^�0M��*l� �}7�)Ƴ:u����T~�B�m_�,�׷iZW�f2nY���#��E�X�U��x{��@��pӲ̱�dyt�I�6���-*$j���>#�"jn���#����Zbs�&�gu}~�3�j�W
ʰ��E4�%�Ζ8���	��y�� jZl���Vg�֠���	�Yх�!ؽ�5ꦀUt���$�I�`]�-�JI�$z�LzN˛ C �1L����4@/��	�VYϞ��y$��� 귀M{��)�% `#�)��1�g�5����M��`^X�N�Q�D^�
��y�M��o��R����{	]�/�����ih�@�Qg��r1�h�O!9�����ݤ�(�K��	rU� ��,Hp�+V�5:߉WU_m_�%����;���A�&޶u+��>Rݫwq�R�w�ލ�ﾋ����L����o���h-õH���ђ�%e��J�g�Bx�\�Jƨ׋�.
�؍E�S j���ڋcA)�9����<ˑ������|/��r'OВ�g�}�x?b]+P!͵�����d:�f�����������]�G��~V_ �lƮ};l�'���:�Ĺ|���~��[��S�×�q$�E�E�����	̐��Ґ����)/��`~�H+�`=��>��C��a��_��Ʀ浆bWW�E�Q7����������?�3��o���>�gf�@�Uo��K�m�(R��m�;lS�,\����7ў)����W.p��[�=����
!�8<ӈ)�g�J3i��������Od^d�x��<��a|����������ŗ^F����(������ã�����_�S��r9��ldu�-�H���%���?��TVj���`L��!�03�"5qV��qj:$L��� ����w<Gm��(�2KBi�%j��je��MN���8{�8A܋k��Ʀ�k,*Gr!E��@�K �ʣ@²h#L2�Ր[7o���k�P��z�t�̬Ր�0}����Dt!F��'���iE�Ҳb�z�672e���Da�LKQ^my����"|����\]���-�c6�fbei'øcm$)z
!?�wn�о���B�u7ÊJ��Q�m[�	���О}hY�
e��\������a9���'pR�&N�w�ov!�E�+���Z�Tj��+�sS�-`"�F=���-Z)&]��(e�
DfqU֫A,�9�He��)2�����	|�'�:����>	v���|�*��N�=(�\,��>��,4���m�d�f�*�I�$�%���9DZ���t��5I�}zz���5	_]��5g�m���}��I�{�o;weӇ^џ��+ʈB�Ke�mw����_� n8�Ӽ8����˧h&*����mJuA+,���E;�:�H�	�TNm�e�g�(@@��,�:�Z�0J�]񐆽�˚���r���zq���m��[~Y�Z>H]f*d��r��)�ONZ�L�<���8s�,yr�z�TjrT>Tl�%�H�+�Aa���eY��~u�I��"�@�y%
	�#L�yd)��s����"OR���r�Mo�����˯`̚� �,�b�Ƶd�*��.�'p��RE*�%7+̣��4QY#7S�c�	��b:��>�,���g1����k�!��]���h�Z��}�	���|/��@�7�����7��?Pf�4�(3RT��e����(?�wddg�/P�>O�]0:�ve�Ni���ˮT�BЪ�Tt��4/P~���#G����p��s��E|�{��'��b4����X���.]a��SӅ('�>����XG��$p�X�c�QdPh���.�=��!�MK�d>f�f��Y��z�n�w��7i��e|�_����Ɵ�~������?�Η,��V�V,ʒMRlBk[�>:ri?��8M���:M�X�AcDZ�D�hc���#5�F�����}��PD@Ǎs���S�j�Z@� Vf��(�[�{��y�����UW�u�\�H-�u��~+�ي�2�J����^Ȥ1rႁ��1i.R%_42As}qV��	�����Jˊ��FKH�bѲ��\/���$�0�,��@�?{���wu�#���d�"�#�C�^�e�cy�=�;��,���ÛՔs��jn��hV�	y2t��d��lX�m��u�ދ�?�68�M�ކ�wߋCo}nx��Ѳr5�(Y�,��m�V6��-|W�O!��%�_�:V\���P%-�vq,���	5O_��]�T��h�S�A�̷��!�8G{��ojb���޺�B��"-� ��ƃ��k��q[���Q
�,�-5���(o̧<M�P�7��X�`'NbE�;B����4�u���4Uu�:݈�m����wU��z�� ��Nw��.��^�3�uy�3���z�[��KJ�Ź�l�h�T���z��G!�U���n\��ݸ���[Y[��J��̟h��h�U$��=��y(���Ԩ�5E�P��Wq�k��z��@�m���eM�Xw��e�:SlV/���j��r�ߧ����T�G���Ӌ7��f��?������ɟ�y|�������?a��F����۱c��6��'rTε���qB�IaV!����:"h�4�&h���*K"�R�"9;Mc��ચ����"��:�,�;�h���Z�{E���̩�D��&���%���j*cj!K�F�H�6�MŰEW�tu(�<X8ކ��S872�iu�F�{+����(���RQ.�~r���@�Q�jNg-<�º�bmq�v��ء'ѕhO��_t{�5��d"��))杴T��B���I�{��Q�˿������ַ�ø<r�	�iZ��{�=�K���P�i�Іx"���sL{���NV˫���2s�x��Y[(T�$&�x_ֿj��`|bS�ҳ�fF�z˭��_�y|�C����e<�ĳ��?�+����s<�سh��7mM_؉լk��o��3* �t��hI����F��0��7���I,3뭉���`Udr��3̛�5�_�����H��@�Uׅ�W���Crq3��QV�*j}� ����I�0��%��~߭zV�L6��5��ˣX����5��Z%s�RS4��ըB�ⵖ��ӪqS덵�S;�#��fݘ�h�yov�O��E����n�c-h����2oN��~T���V+ϩ����c�����`�-�Xi���ņ�7b�u�бi+��:0E�n��r"�n�
�A���&-���L���9计���Ǟ@&�D��4iu�!
9/�#�u+o.r&����X�6g]����LEaz�mAA+���V���b��j�\
��m��}��p��7��+fK��)�)�5Y5�<��&uԥi���F=�Yr��N���DXG�F��h��Dt-�j,�.LP4��y�՛���4V!����Հ��^�w��&��������:0n�%'P"x�vn[�O|��x��wc��Z�ݦ�D�ku��I3�R��۵dݱZ�_a�a�JZnxg�'	�c�T2U]O:�|�ɺU��ZZ,����� kO�9G�1ǹ������G�6�9����:��������᳟�,>A |��	�aVP��^�G,��55F@�x���"���5߯9���	runJ9�\P%�yaj^���Db����S�&g2�^hey��H��Ӣ���|/���FY��q�Z��l�$ݓ�����%�n^���+�l&�{�-R��#�5��K�g�7h$_����M!�T�h B��F��^*��l[}_yY`y5�QѤ�Ŧ�rn���]�Gr�׹-��h�j�{��TO��ajj
�Ϝ2`?�K4G�_�$[$2yDc�v���38s���K����i�6H��3�J�.�PH9Q�4Oy�sƦE���
�H0l��I�ieh�Jk�X����N�:2���Ъ>Di���D�|>�wb�ڵ���F�_,㟾�������#H&	"̳�ITf�d��/��JE��
c�Hx
Uc?�����4	�Z��Kd-26K�l:��Ye�Ty�a����G&ԥ�(Z�L���upuv�E(`}$�f2��~TnR��K��w��g�-]�I�0��ի?��^z��r�L�?�����*�I
=:�`!�^%'O�&̏M��<��c����eJ���z�A�$#�۾w�u-��;�}�:�jЊS�	j�qD�j�Z0Ǻ��m�ns�֜�H���VD[��ѿ
52A��lx�Q%��]#���dLV#���@�	A�'�T���\���0�*#Q�b�Ԍ���u�rU�Qv����d�j�xR���a�86�b���Z��Wx�-7���j��.*a
���/����9���,"�ϒ	>�?�ʈ�	��2.�z	E�`�`�k��s�L:���;V�]o������9
�l��D1Z��5fV�����r��rH�+��&�J�jΖ�b.D*v��Q�},��%��<�R�	�~KY2���%蝬��%)��4TJ�S`\yZ�+N+d��Jd��BQ�6��j�S��w#�h���>t~ԥ�Qغh�5���"O�X��՝��߆_��P��zIN�-B��T�߽D+�CaK��
ZVH�i�$~�Z���2�'��|�	Q_y�V�,�J�tB��d=�Q&i�����6߬N�J5�#-h��޽��aZr'��v۝�S�p����W��������7߇�Hgs6DQ�7�EV��0ϝ;m������j3i�mF����Jvm��۶1OՌ«�(e'm��
���$��Q]�""�Z�5�S!G�r���Zp��$f�ճ��9K�Dœ�I���@\cQA׶m�&��E9���I��<�@Y<QJ�g�@�:�M�Z��򤧤�ؖ�by�;{�,^8|i�a:�f�����ZD�M�%MP�o���jLN���ŋ��![
��)��*i<Ԕ/�[4(�g�����$C�:�%�.�|��{�b����@��ּ��`�:����C-,��Y�2͓��z�|��L�R���(�f��I�'R�_�h]��dt� ��5w��H^H��
����/�
�Q�c�A��w��;n���>VB�'�̳����i�P�"�j!U��D�UA&+^��[X=�J�"~��~������6�Z�)ScS�؞e�I���Dך�p�t`>M!D��R�1�kN�}
�t����Q�.
�>WȲ��25�Z[6nb����Y%q��9K����_Ha��E���n�a�������c��Z�7��:i����Ǎ7��>�I�߸�\{+Vm%17#C@MtΞǹ���&h�=�](c>��@k��v�%3���ͩ۫*�u�SI��J"*���٪[R��
_�sK�t�%3QX��d��"R`�?j�Dx	kѯ4m[Y��h�S�����l%<*�}�$��GnZ��Zv����}
P
1���hE�,R�9��M`ݚA��ށm4�lyen̊d�P3e��� ���e�j������F=6�RZ�4S�����L��z�&��٫���Mٱ����#�Q�����^�5�ic-*�r2����&Q_U�K#�
�1a�0�Z�UKj�ܺ��;������Dcmʉr��϶P@n9l�m-=�>%���D� ���Hőr�F~Z"px���&�3��|��D�|~�����h��l ˗6޹s'z��p���h�|�~��;��{��DgG'��M�Xm)�!"k��c�yԒOᐗ���:i���hz�\?*�Hz̏^�+�>�ً�(IHO�"��Dvn��58?e�����H>�i�9Om]+�?��B<h�g6�^K��M��e��6VZ�P�����*����={�"�h��0�7�YW�u�/�&�6]���!*��H��O=*�$yT�B�se�F�غy�-ԟ�H��S����0?�z�1�tћ�B�.E�Q��<A�H�딦�i,[c�/=��/~	s杙'�$|S3sl�ÔIՎ%+�I�5g2�<�+EEjF�
M4J#�5����SzgSX�W��2A�F ���r��װvM/�z���ԧ>�O|�'q��v
*��Ԑ�w~��)���45=�g������F�7�F���,�����d3�f�-��U;��+���������bՁެ،k��@ۊ��X���49[cJ)�Q5'EK{�h]���#�E�ZY�Z���m9	j���Ͱ�i�%�d�4�O�Éï"=��M��������M[�G�2@m�E�brl�G.arb�£�XK7*�0v�w���\���5\����Fp��N�I6ad"��t��pGۙO��g�k��l*�k�X��P�~XIZym��l���Q��"bu'i�1����1��J&�Ԛ�?Z��t	��y
�&�̤�Ȑ
�M6���,6	��JQs̨�8����{p��{�9*�W��72KeL�37���O����,9KQ�r1�q��qk ������o�tM�B�3G�!=�� �7��?T�j?��rR^{}� �M_���<���=:�t]�+���w݇�ﾑ�V
�� Nʆ$�����=�X�u�Y[|�`'�Tw���T�.y&�"1��<�\j��KL�Z��ܤъ�����[/o���2�By��3��|���2���+��~���q�Fdh}iޜ���Pu�d���j��-!�/h��T���2�K�`aj��<=�iSK'��6&(�IyT��
i
{ғGV�R3��V�ba��w���DX����U+��'�i��x��F����OY�h��řE
��>x�Ȭ���t��Bok1�>�UC"��0"�y�j�PXsQ�i�۶;7��B�� W%x����r���� 8�Mgf&1;=e
��B�Q�3�c�鷎��R��!+K�@:o�"�ٶm�f%ZZZ��tX n�Gত�5O��iq���X�'1otJZV�i|\�e$1<�����{r���k�8�P�eʌÄ̰\�4�\Ӟg�R�����O}�6��֍U�h���cL�Ѫ��jǞ=;���� ��O�c�~��>���}��o~
��K�43W%_�4�uy�f쭌�HD``�jw�Sg~��г��lo'_���$@*�$��+��R�XA��_��x���[�,�Ә�������f��\I߹r2�*-�%Vt��v��ORk��y.
9�I�MK���X��Gbrs��I�q�ڸ��H/&QHi��<�/^&�i���˃���KgiT�ct��ǟ=�����[H�1$uL�f13ZL̥H�m+��!��YMAC���}ms�m�am���9�M�n)���Z��bs�q� @�i���wK��<���3>�.AuM���xB��/ˋM.���j"-�i��v��/`f�"5X͓��N�rT�Y�tK,���r��ضZ�N��Ȉ�5'0ȩ�P�d�P�y�1�YI�.�5�ԃ�]�9���D�-��U2��8Q�������?ߣ��UWk�:�$A� ��]�=k3l�������e����xw#5���g��,;�$�%%��$˃s�?���ĭ���[Lxj�4�kF�秵⬭GB&�Qxi�
*�T��1�S�����۶�����o������k9ģ~���&w����0��q2�		�W��׿�o8y�4y���'O�s���MF��_DoO�y�YsZ]�!Z����&�������1������<��itt�w�	?����/�}(�&�������+���1͵���%+��`�q�%u�F�m��4m�M��5�I�@�Y݊��'�7p�=M�����Q��M�a�w�t-���Ff�<f.���ql_ۇ�vl��thU�S�/�i�i9��r�#�xph�v�=�ܸL�����"�ʓ���6Sω"�T��	��^�O����}���^�5�}��X������T�/���^>������G��vT/��<*�P�O�[��m�x�J^@�O�fkIR�h-+H
��D��l�u�[�:{�Pǚ�c�λ�3҄|,��@ B��֑���G�,���v�tw����\�o��x��o��+�1@��*r���0�U+�J�C5�����ə�B�����:���ּ��������,M���J���JT@����D�Zy	�׬�,��@��҆�|�;�Sh�k����	���0QzÈ�#h���`��-�ƆG����=n�}�0�H�/�����|�^����al*����Y9q	��Z��OS��ރt�N�#�4��b�n:;py.b:ˠ�J`]�^_�D�ucӡY�Wȥ��V����~ܦ+W@wy/"�<*V5V�43fgH������g�K@{��ޣ|F(���;G��\М,2��V�� ۙwkGk>��c���d�%̳N��bk�9�U82��$)bRc�˂63��RsG������P��@Z��6���Wo��^�m�̼dT�NW��U������������W��1�.�w���)�D<�٩�ޞv|�#?�m[7�}h=S��֘���'+���*�Y
)Mё�N��:��&�/-Q����]��������YLg{��,3�z["o�_<,5�ak�z���I�9[�i��W��<�;������/1%��T*��_Z��C PLQ�(h!`,�js�g�*����~���������}Ϊ$�;������d�
�m��K�v5F(��샛|����j���U�s�)�;���JX*�	8E���U�e�X�'k�"�6�ć~�~��ͷ���xۛ�]�ߌ�k:�-�j_Bza/<�$r�9~�
G~,�'��عe�K��4e�K���B���n\MKY��A� ��m�Q4�D�%�At*Zh����S�����Yh�D���a��Ӧ�]Z@8M��jz6�`R;5���7����;�i1ZkQ�>����[��F��6_�,��慉�t�V�E(Vp6�&D�<�\��zG^<��3#8��y�r��r�ځ�Ib���������sGy�Y��H	/>��-Q�n�JStsgj�LP=�Od�B������r�j3"�N]Cb>F��U#b&���Fm�<�,���s�<-5_[;w�Esg?��jUK�ȳ�fݕ�MQ��J#��{|����"���g�$���gM��Q�j*e���J�"�u��چ�e�y����;�m��Ԥy���2\`������19���b�\3��~�{��'1�t��Ԁ.�����ZL��tݍ��[бi���%
ry7j9FY'�R�`ҟ.�yM����f��ݡ���i�������ˉ��-���m��L�����j����!��-�b���`���n�C�B����U��bm_��#��L��Am�a�u�n���pX�
�=;���ۮC<!��	�������X��s��2�4��(��&�Spa�al��t�%K`]���Q�)X�Ii�Z ��"J!Qִ�W�3_��Z][k�nt��S��n�
4m�5���F՗4�F�4�M9�4�۞]N?jӳ�$��_�1�`��o�X^�*���t9I�V^�W����.l\ۋ;n9�
T�I�ŭ���@������"-�,�
; ���RsS����!�s�	��r����'R��J���V����h�)��ܬy�J9���$_�Y�4�@!�Α?�4��h4��$ﴚ�V�_�f�v�eE-���~�5�G��@Cx�=q/�]_��遴ɇ�}%W��rRu�X�(2*���M>����U�O��Y�������"\�-�
B��z��Uf�l
T�gfR���i�5����������>�_���q;u�Y��y*!ʬ%�z��j.9�J~x����"F9\&�hb���]��-�Ju=gWZ��<-�h7^��
g���uƦ�>�Y�1��5);�1��TlՓ���I�
0�5�G�4'E�h�ug3L�;�M�X�%͍��V�;�S
�x����bQMYѸ��]ئ,�}�3�y@���)�ʹq??��'�x[�E��!Q��4r�.��z�i<���0|nc38u�~����w���0~�	|��'��G�ԓ���c/���W)�XA����B���L���Xh1M�U�Z��C��ʭB%b_��xв;%Z�>S���e��0�Xf�Ld�c�]z�	�AB��C��^1P.������h�B��*�<�.��rވ�RSTv��o`��/^F.�F@Pt�:���n��F�Z&�]�on8t�P����5��
˭��p�ց�6����7�y�$�˲z�,�˼�4Ἐ�&H�ɓ�h!�׮���C@gf��Lq�,��լ���^��&A��%���H3^
�&9�6K�s��m�;��k���I]Y|�R�%�c�@���x��W�Xj��W�I��Ѭ5���c�Da�Vt#JEb��q
A�N����V��D�w���I��h�Cٜ.�G�%cXN��ZU�>����WhO�m��H)��:V٭0vM�(��I�R�fݠ����I�T>ĀdV)ez��λ�^usJh�cvM�b^ ���
�o�P�ؽ�e�y�Gl����i{�����qJ�\��N���sv��?�����D�S06������QpG�(���5���u�[�b�X@A��U���������u�Њ���f�:z�rf��G��DlY,9r�N�bRB��Vv��eU�V��ʕ�X9��mq�_�X�<;;;x�.���a�M����C�P�`ph��ן:�{�!����n�@O�ь����R������c�˰��ɍ_��4��zS� �bL�2E���iCcVʹh����um��5�WNR�%@kE���.��<T�p��k	+a�[[�b�es$1֋ϳ�|.mQ��B|���ox�#�.j��U��O��u)/�E�,&������sG���h=��
���|3��@�޻n���Ο>�B�J�&^�^ծ�;S8h��Z���&�۾A?Z�ơ+Ym�Ӌ|:g��}��8�.m��s�1�a�!'2���L�[�v5��ߎ\͍'_���	*T0�cܥ�b�o����|@L'x��(N���7܅H<�YZ
�L��A)�8+h��m����q���������jZ��k֯�ν{p��w�����JXXLP�3�9"PP˲�i�ǌ�F�};���5�Xe�xl���I�h�<)5Y�Lb̑r<]�nC��������+I�$6j���km�,��\r�X�݊�5�Ě>,�WW�־�hcŊ~��4.���	��-gy�ɽ���xL�@昲رk�E���#py���C��"�[hAR�Dh��	����|źY
�O�TV��O���F�����[�@�ƭ�'`�h��yY?�Z��+u�HV!ږ+�����KMQFDS��H�����l��k$]�ll�-o<acA�˺O�Y�e�]��~�=}� )�-.�.��WQ�(���ن��󘟾ĳl���\�P��\���j�{��V
��lk���@�UFˇ��oy��qcP�O��;ʗ3^�P��i�z�Q>]���Q��\u����h�`�.?i̬�L�:5OI�Qyб�u	��RW�,=ǻ����'�u�T[8���ϫ7��Ο6}O`��ѽ�yu7��/7�'ek����>e�Vټm�ͣ:y������G^���f@�v���V�u��n�M׬D��M��2���a�>u��e�-زa%.\8�:hƍ7ހM��`��m.l+�W�\i��\{-nP\�}{q݁p�^w-n���۷{��Î;�e�flذ�W�!N^��u���[�s�سصc���]Ÿ06��?��8����mEؙͭ�	ʤ�' y������dqHբI������}ذ�ˬ���������\>d��i��2�T���F������o��c����n$%�Cr�r���S�ۿ�
���GL���`~�������a�d_���}3�	6+��(���#�ei]���"��%��_�R ��hЇ"�{R]�^�F�T�Km����7~_�5�zӰC�x#�UO���S��M�mX�]����x�Ջ�<�)^�C�V�3�<���,��TGN��ԅ9����:066B�����c%�����֛q`�j�]�a�"4yw�݅C7_��o܋]{�`��5���҆����n��}x������?��&#��Յ�m��ɬ����H&���^��+��[c�
QT�2��`1S1�W�:����옕��z"��CW"�1�'�O�Hd��P�V�x%��i�`��'�h6��@?���҉�VP������&�j�"��P(xY�LIH���I`#�S���_��"0�(`j6��E-?Ta�U,:��_�4 �*M���ˡ�o��k`��F���I�O�E����1%;�L���[H\ګ>�^�u�PoԽx����oӣ?��� �ږ�n���up�}cj�'��a!C˚V�ޯ8����hrZ�'gR%�K�^����0Y�rS�,5W	+H{���q����Nk9��J��M�M)\u�*S��Y�u@K��z`�xM����ҩ��aJ�뀡��kN��\J��o��� z�ڄ��I;�;mLJ��P��!�#��kB~���ك��>����kS=�߶��i��{t͒#xIۿx�t��"�t[1�R(�r(`5y��[�x��1,.,�����7�c!�R�\���EQ�x�\�s-b�V4�O�)�_>�'��=M��t�)L��L�p��!ʥ�)���WMQލO�����בr٪��OY�#'ȯ�-��e*Y�}$�_đ��`�����y�U�l&�gS)v�Pq��$�F;�L�U�y���`G%_�ֲvH�j�#鴜�u{�`UXeFK�33���Hf��;-)�������z)��8~LV�-����Q��V)fϾp
��/�_���7�+�5�Ɣ3�2���8q������?I�5��|��
�B���N/o;�n����Syq�-<M�צ�S8Y���/O���k�~��!�pc�PllW����uViS]�E*�_���E %������q��$�����\��װ�V�=$E�Ī�
��@��h�ʆ��KO�����=kI0~$X���j?�<!T�HK�K(өL.�C8�L���L�i��R4Ȩɳ"4��XQ̃9���_��7G���v?�I�|}U��M�iY�*��=Y�cն�L;���B��F�Z��Q���Ej_�S�8y�"�y�0^z�%d�IDC~F�p3V����-l��C\ك����7@OoZ7�:˺Vh0��DS|z1M�dc$�i�n*WB��"@.Y�;��P%�j�S����`h�.��w-�Z�}1g��\c����)�(�5N�~oKlwY�)Y��V_<`S\��o����׽�6�vG���� =h<%����&��vF�GH3 Y35�O{gAd	�H���E�#�V�d4�`IqMo�����h�.�V��~�������F�ըo��y���\J�"+�P9��) S7�7�]�ޞ#3ʩCA��}E�X ب���I����SL[ǲ�����է�,1��m����1���������)/na3�d��>�O�u���G?����%�S�hfj��7'��@RcR��C�e�D���ް9{�����l�<b%��k�.ֳ�</e��Ri��5k��
��fS����G*���&5F�UM��2�L ���ے�|�>����KY���20�؊�*:wRZ}�ޖ8
�]vPlR
��
��DL<�'�+"�z��I�!�#�EO^�aʠ��<b�s(�S�ˢ����Gu�G	r(�Bx��s��/�)~�3��/��_���o_����9��?<���7_�K'��u��J.O�2�Jq�@�����O_�����;�������;��ZTςH͗��]��5A;����ۚ�� 58[��Լ�uy�g��,�2]�~�f︊��^񀆠H����|OY���T��VS�o��]瘀gcd(!��e��UH?�bt��FZM�c�;{�"��ￌ����_����=���_��K8|z�&�"��_��v��H0
ۣ�	E���J��f�\n���Gc��J�#6��Rw9o�_{�֝mvB@K!�k�_�_|�t�eg�zw�CώkQ�aBV	7O�WW��X�{�Ti�9�o~�a<��QLN-���>{	Sc��σ;�	o�[pݡk��1�(���T	M$�����?�g.�8���\ro�4����*�
ZK~$k�+6`p��(��NP3����r�*�(��J�9��Ķ�qg�jcGJ����HL�^����k����*[�kO(/�[D�������I�5&!gj��E������=�:ڢ�r������{$ )x����Kصk�|�m˖i�:F�AᇭՕV� ɒ�����iV��g4�nݡʳ��oi�o�D��0�sNȫ���姐M���"!� [�����G���m ��ʓ X<+��^m��>r����2�|������h3��
�������팃�SY�z����m��f6���l?��v��Hc�b��e���T��$��.�|�I�ɇ�,���~��L�PI��BT ����̌�Hk�H�?��@��QD�_H&���q3�3�b��ϝ;g֧jD�x�M�]`٧g�i�kNJ��V���r�u�˼�J����¨5iI��,73�O�d�H/�4S�e��0K���]���TR@��:aV	�RRY��3���\�%�,X@��FBz���������y�Y�ޟ�/����	>�ſ��/�&�F�H�w*��2��)�T!H_���Z���BhA"�D��R��W�o˥�/AQa�� ��5�y�̣��
Q�5��m^��&��������F��A��1�e�R���@�#�j�e�d����_�O��JD9\�`��jQ(��W�~�\G[�M~ڴc��.	856����_���P��rn���"�҇HO+fɵh>թ�߳�rЌ�)������8rv/�r�>�'�{���%�9q�����
1CM�'�R`7S��uG�I+(�>�Ǧ�kP�t�*�L�d�ݫ"�_��՛�K�����$�l��$���#WvH�*�øˉ'Lp�"��"�d�b.j���p��|_�L@ˉH�g>~�N�A���.�F���%S-�*n>xV�\�L&�ɉ1l۲���E�e;qJ!}�c!]`�Ȥ�Xpnx�'fh�(���0OfJ��`�����D��߆�����}�t��D2g��B��K!�i��$|�t����v�G�ĝ"騫Z]�U֡��&#B��%�78G��Wt�|�~X�q4
I���S�<�J�!O��~�8�
N�:��`��Y�/f�
���X�y���@k��|�q�XV/B�5EPi�P8��3?�^�_�M!J�Bz����#�b��pX�.G�v�ʢ?1����;���Y�O	w2�����ٜ�;ev�k��e�eYN�R�$[P��d*i�G�,�ի(H �Ik��';�>�ҭʲ�uե�N�Q�%/%�(AP������r;��c�������mw9�f�UL缓��؈=YzƂ̳�}r@`���2�}��Is���cl�:��rbM(����s�
*vo[�֐��ha
��D
>��*���>�ݻ=���^�ˇ�`fzs�sX\L��w��es����SV?��f���~ZMatt��cxxc�c������Q�Њٲ}'�?x�1�F{��wZ�j[����K����A��Uw*��\�R�X&�w�v����<>�
sU�x[��헚č��`�`�͇����q��Yޣ��ⷉ��n�A��Qd���(׼! ؊�p��=4[�L�k��� <�����)U�����%�"jeʉ
�m�ԺqUw���R�a#+���c���<��"fh1g3����,���ޙ��Q���4�����쬆+Jv�2E�/	ܮ(j<vbh��eye�����5��Z�`[�5�Q��P���3؅�7B{w���|�"�g
�ϋ(���������̧�ŵ�vr���\Z�/J��cV˹W���].�0������
��cO�����c>
)O3���#pqn����݇��G���O<��Q���\NKdy(��h�ֵ4�5���)c9U�#t����;�iGl�2�-�P�ʪ6�U�o�ca�{��寰��eVm@����M6����h�6#-��s�`���46�T2M��3f�(�!���\k� &gs��x��E�N$i�ɚ�S��U�u$b��W��K�"�a7	�Dm��D��cW��9�5��O{72d��FM��}������D�����tM �#&����	��b���紇��9�眳5ZL[�Ư��Cޯ6�?k�J	1��VDp��a�==EЦFZ�^y��5#�f�즵<����H[���X�ɭK(���,n�� ���7�Q��H�
m�z�E���n�U��+'�
�C��ގ���䅦c~St�Z�e|m�.H���B\.&��H��c�j�;��vuuY���@@kz?�%kV��E�`$BGG+�P��Y� B����_�<:gʍ�w@�*��p~뚝�fW���c}�5��K)���;����m��U�5�Mݰ>����h!}��b~!E�� �+�WZM�"g��������؈[�C�ġ��յ��S��'�E87塧��Vt�̧�y�>�8��<���	�8�_���g��t�E
�EZy��L�������g,"�ٳgq��I<��x��gq��I[ht�5�F���+x���M>�v?�1����0���G�_���A0jcY�*>����=���N}�F5
n5ĲzvQ*y�r�� ���Y�T��������PB���E`�N��\T��0i�f���IK+5)��6��I</�f�A3g�Zy���E�s�a�NkI�"ȁP�ظ�D��xh�֯]��)���[ �N�^~�KN4R��@"�$݈~X`�Z�~����A���&p����N�<��G-��۷�{�ĤY~/�,�k)���x��رWF��si�pbc�y>�C,�Á�k�1���@F���3�p��,_Њ0�q�����(#�KP�b5�B!��~'O�f��)@|&Di^���K��fh�yO�#K]�<y� GAJae��n�h<�-[���x�,���5���^��՚U�<��z�B����lբ��*+Y���WmV����.^9��[e�t��݁	�Z�#1C+��Y%��~� ��Y\�Z���W��W^���ØI���x��N���[�WG6��Q���w��ؕ��<��b�@a �_][�ǃ�<�x���څ��{�rﵨ�Z1���y��KP];xW�8�:��Mt����*��1)6�Vh�#�����J���e{حN{��n<oG�o��߰��?֓��f
�0��[/`��8���g�-(*��x�ﭠ�=��0i�f�E�Cd�%~S�C�]�;Xt|��ĚU=(j�VIݜ��Ɍb`1��S*J��e`���"��d���^_n0� H�尿�Bj��v�9�C g�L��VA:��yK�4�FÈ�CԄ�1>6��^z�{�a|�[���>d�=�y���G��O��1	��T4�L�<*"��#~Z��g2���{hQh�C��������<7���I�i|�6�K�	��W;�Vv�h��� �=	�X<����;w#����*�HRH��QW�ާ�����p��>�)�j��/��x��1�X9�iZh��(���Sgαb|���e�&b�ꦙ`���i�y+��Ri��Z�c�@�9�rt�孶��b�P��{����7��-�����k�X��|��y��#Ô���<q
� 늆�N4K�a5\�2�3��?���_B���C��bϖN4�ME�=�F�3(�h�uZpK;o�+7yd��N�&5�"`	Ju΀MV��@ֱ��kZIʛ����dx�йOJ�<�]�p��y����{��/Z7�/�ʶ�B���3U�� ��O�1��gz��խ��c�? #K��^�:whd`rN�3�;�s ��%R%Q���mٖi[ג(ɔ�������,��}J��3w����ĝ�� ��������f8+��-L�9}N�
_}������qz�2��'��o޹r�`۾+{s�;z� d)�F�nT���� ���)�R�����Ħq�]*��`/�����L�Ayz���6./��G� \�SIǵI!<�iHz��9Iϒe��v��ۍ7ݨ��Y-X&޲�}�E[�ٻal��p�
K� ���P���g\7� �
�9�蟞�0
��� �9��F�\H}��T<�{$��YK�*D���Ԑ��ö��Gl��{|�.�X�.ɲR��N�'m��|к����ٲ��X�����r䒽���� KnEL����^�L=�q뎐PV��HU�*�����͘ʈY3-k`����w�Yv���7$|��+��E!+8���G�w�*H�ǃupv��Q�	�$��<�3]�Y��zƨAײ���ʊ4���ѐ�k5�R�|*Ҷ��gl8o���]�h	e6�G�)�I����:�˙���~ߵ�m�|0�&Bc<��������x۲da�B��;v,���Y\=X�Bl�%���"h�.�bخ����������d�����_���mߐP;"+��Q�<���9r�O�Y��>�E��O}�~�7����o�#��_����?����B�ᨦ�A�����#|�Pa+'\��r�㕺E���s��y���HX��(Ĩ��c8�6�@�!2���[o���:��С�
��zO�q�&mΕ�%Eѿp�CH���-�e��[R����ܴ�6l�"���c�6mۦg�%Ҳ��"efU�\��9+���s/����o>��=�����	q�GFmD��L*
��VQ^�.j�\�&Xo&J�N�l	�ji��	ŕ3E������z�p��lHA�[���k�VZZ������a$��b��%!���[+=$��o����$�}��h]�rU��h�u�!��p�)v��?�W�c�9x[���i*��[O+B3����c����ͥ��E���d33�~�˲��,���Qxٚx�pJ,Y@h���j(V�
7���Q����0�k�W��p��2�0i˵;vv����|�\~���O�,^"�<�w�,��
�L4�5�� @"�z�0R�>;yꂝ8}I��k���Q�������?d�x�����~����G��?�����i�xǃ"x �f/N�Q1�TWZ��� �^��0M���$��w�h�h��	�����-^o_���[vv�fkc�m�#�������t���cVh�l��g���-).�ҶR���˒Hؙ3���R���:�gvU�]��ݯ��Aa��{��Jʫ�MV�K	���gl���]��m��.�fl��)�,9�.-�!)m�;�8����;����P��^�?�;���!�<�w7W�We���D<���MAj�Ną�/Fǘ�����#���w�w���bv�{md(-�ڶj��fg��tEx!�O�݊�J�$� 1:��0yŅ]�.�3�?/0�e.�-�s�ؙA���������~�W~�>�Ϩ��D�E�X�('�'|�qY'c�c6::n#��ҔR��*���m�O��?��O���������ǟrW:��ȑ*�j�]�aD7xG_�_Od܄�t�?�e<�*�A��9<$'�|����o�|>#�A�/V��l/����cꗪ���p��f������"5Z)�����e����3va~Զ�3���qfƎ�qJJ�vFi��O�������]�4#��.β���-�T*�-7�"~�v���S��P�P����xjL��%zXC��5�}Ĭ� �$6�6�HM����z���s_��-�MK�yٖ�ӂUK��Go�U)�>KȺ[��I�fI��)��sylW���.�)h��9��Bl3�<r/�x�3�cM�/W&��:�0�Q��ʲ �0V|�VB��|�'�
�ܥ	�!D��89��~��]7��@�xE��ҽ'��u�1�m\�hJ��UN��c5�ʩ9Z�)A�2�f����\�
?Y#D�0�ŅE�-�pW���3q�������;O���펻����h��?f��������A��?�C���$�D����ܢ��g�TH��!��|lj%�U���@�O0�(�U�J&���.��9�����X�*x]"�E��z�"a}) ��zV�pKٌ��(9t�z����{?j=�m�gܖZCV��fr�͕36�"����DjBVˠ5VVmĬ�*k���R�ci�u!�R�lS�s6-�xa�$�������v���v�O���eW���+;�$"l���Y	8Y�u1u~[�	HQ�A�( �(�۸�~��]W�:ߡxMP�jV���"OMyѢn�\��o��C��U�Yy/׮68<��ȑ�i�8�mp�	�֨��}Sb�V��",�ݷ���-b�"Z	M\���Dyv����[�I��]�T�IHI\��'��8�
n�(0+4+Ӂ��.����c'~�$��k�������O��}�_Q�;�y�f۰a�� �U��8������8��fP|:bp���G^�D���Nn�l�3s�����_����OvF�S)�h>�	��/T�� �<E����\��{o��B�H�m���l=�1�-�?3�Y�t�}wJkgUB�wé�b�',T���;��nU�I�(����#�&&'}|�i�{��o��7qHˊdb
-ne�c��B-��6_7dc�rj�����������ə��$�T@�ND!�$ؔ\��lᡌ�����X��cMi��E[S����Ƣ�-[�V���j��ʜ�d�ҢMժ�E;|����p?|[=�����'��c�X�ϡ�
�Y��\�YFx���z;�����q?��d��bMK�9V�j�Ԛ�%�,ωJ7�Kؠ`�핰��儬����#�	}����W�NU��lgOu��R}��YY�����9�1�`Ir�\P�R�(fx�%'�Wp#p�����#X��Be����|�-���������aN���*�����8�Ge��~��7U;Z��1\��Y|�5�'eSK�I�U;��E+J㉧��49��W���Sg�r���?����o���v┏1�G�i�F�Ѻ�1}ڼ~�t�ˣ�b}�� �^\��$C�	��� <L�i
�2�/U�V����h���z�6|���j��b��$��VӶ(A7S�v���ʃ8]iؔp^� F��6�ա�B���I�y��v��?hw��Gl�}o����v�=&��J�f$�41�w�"�x}/���u��V�qn�͛�WB|�!���������Y}̚c?T��He5^�Z�&������W����4R\���Va{$�c�>l;��Y�ZC�q~�Kvw�pͳ�	�	����ܥ"3�t�,I�0��.�(8t�5�ݢQz4ى�	�1���/�忲_���ge�+mZ�K�{�a�=�
�&�0U|y�`����}����cGO�K����T��Z3j�_)VM�-�`�F��2c����Nq�}�>���G���+��|�=�k�6��C�mK���
�����]R�ap�r��a���ʉ,"߻s�=x�=��~����w���{l��=C�6��Y��q�)������K�z����1�������n��6�2�q)����{{�lDߏ*�֭&���Kଭ�k�*KSVY��եik.N���%]g��0k�D�W���w�Y��{qn�� |j� Ex�#A�Ϛ�{��Ν���%j6�^����������U�O���9	��m�ې����X�r�*gl��Q	�9	�UP�i,���u��{���K�+��^�`n*Jh��s�~�Zܥ�YW��|���Q$4Úm���I�߷�v��n�Y
�'SЅ,<}�{�
txs^8���;4��ÂljT%܅�C�}64�/܇2���|��I)#m�Ԍ����F�,��@uݲ�f��4A���sO�� L��e�o������?�������?�o>�q~֦f����i�Ɠ/٧?������G������?���Y+V��x� ��=66&�$�3�(�EDD�����@Sx��>�?i�Ø����X��c"����$�x�lY�YqM}~Ĳ;v�Y�7��=v���������x����b��n���v+e7ق�����'�V����d�!]S;o���?j{�����ڡw�6���ٴ��{��\�i�`�b`u,��RC�����p��D�������\f��Ҭ�«������y�x�qv\�>3bǆmP�|yi�����\�ZW�.�l�=���"����V)V�Bb����υ��+�cr<G�1^������Jx���5�7��I`̬T.�9kL�a��O�����?�W_yնn٦�b�*+��B��(Fe���=��v�*�>��+��z���Lf�+_��}��?v��OXE̂2c�wf�a5�(�n���ZW�w�k>P�)�wc���n�-�'m���^C�8S�����L�,�N0�>1._|/F��f�y��Q0�ob62���['l��Q�2>�{��I�Qd��~	�q1�Q��9�*h�`�V4�v�m߾�~�{�-o����9���p�a���%s#~�ɂi�#���%��R���,Z��Z�V�D��{~,�(H��RL�Y{XV}׬�/�Vn��tL��������l�Ě�}��h[��qD�m�w�F2eΖm����e����e����֣�S%�<д�\Æ�*�5g��Yk.�U=��\�`�6��P�l��,�yKՖ��#�ZE�<����6����n�nW���b��Ey�]1�����-�6[~���Zͯ-�_��ٕʷWT��r\��e�.v�|=��O�YU�Ř�P�����,��J�:�����c�P��W)2!��,c���_�$��Z�^>9�g��m����L�3�����H�WV�W��J{�:w�^z�9{������/�׾����|ɾ��'�g^�j#i�mE�H2�z8-\W[mYJ��6�v�ݼW���q14_������,��AA����nd)Nj[E|`�)k�d�oF`��NX����}yP_W��L�A��r�k�갎�L�`0@�Nbh��7l�-�n��}7���ֿe���<`ɉ-���ַs���Ɇ���m۝�َ;�ͷ�i���[��������"�J5+0�4�n	b=hL�`U&� ����~�~�>�E�N#B̤qV��#!�N����K�������B�
f�Sꩨ�<C��� F��bZy{�����ZovDP��Q�w�\o��{�j�Y��ЧʡS�l�iw�q���&i�	��j�J�g���a���_3�M��S.h�^?�`�N|��k�� ]�9#| �"W324�����]���w���l��m�g�^�+
8�k�
0n�{6l�n�Q������u
��P���O��Ý�x ������'�رcBɜKCgb�(�:��K��uu @����y�g�z�Q�g������+~�@N0�W���J�ۑ#�lna�u��r��ݲ;o���񶻐��-���o�bO=��m߱SV`�|�n۹m��n����s3���S��@�]\.zrj3;򻂣�X�����q�Gm���;|Ӎ�c�<���W^�0��w�}�+gx"�7��?��g�S��}��q���;ݸ��1����P��Zu��[l��-�=����Wv�ڪ6�e?��G����倄߀m��o�}��������}���G�a��#��]��[���7����a�����~��#��f�총Flb0c��n�����{�������m��vж���@����jo�n����}�G?d�<�r7H9��U�'�z���|�=0�>1>:�B��SV�b-@�sE��;��2J)\�C����u�~'�'}Ґo(!�n�DO�m�p�m�c��OH�R����xᤝ�TR)Y�	{讽61 ��+��l�hV$-^91c'�I�o�f$�Ϋ���*>���S�1]��م��ΗmiY�d�O��b�a�5c2o��|<��>�g��>��!>����{,�'��UNo`H�*|w�WSC9�|�ʲ��L�V�.��*�,bt����#'�3���z$b�>��+�0�������+m4hY���[vt��o�bٍ�]��Y<)�7�e�%�7Y#5`�L�V$�[1[l+*����nV�����q)6��N0i��s�k��51�.��%B(����K\D��
�֪l-	<�
g$�V�WfxF��n��w�oW�/��JQ�*�݇Gle�jǏL[òV���fx���֪,���/�W}솶"� p�����z�i��	����ǘS���4u��D4�!ă�!D5|�	}���4��I��pF08��6�4%!�J���co�g?�Y;q�mݺU0�?��)y֑6�OܲQ�=Q�Fp� �w���4�\-)B�}��P߈��fge�l�՜�So���9w���Sl��k��:R6Ȕ�a�xF����jB�]��fҹb!���?+s�Ϝ��ٹ����K�W�k�e7ݰ�~��KJ1�����^����.�?/Kq���a)�^����v��q;s��M�M����볿o�6m�l����1��'>�M}�rܣl}�=��ƍc��^�	�_��W$�mӦ�vםw0ܬ�1�ڰ��/��>�eK�v���Մ5Y4,M`��� ���/8;��!���fJV�rq�]��o���>9?�g��ﱛo�c��)_��i<秃��1n��G�no�M?�VҶl�}�����;w�{�ض�C6�OضMy��a���nط�Ǻ��d�&���m�8,+y�ؽ���f������.���"`����q�����~�R@ţ%Pfp��]?�I��#���э/�)X^�
t�DwE*�,a�!�t�obZ����X��_d������-�<dť���0c�>r�.�וw��31	�}6��Sү�H
9�ʀ�Tڪ �d-�F%��'�q"4Q��R�f��&���Xf�&뛸�6ܠ�6��jܦW������LM���o(�¾v�RIy
��'�g��)J��oH#Ă	*i[�)@���?O���'�紅�)[�����U� 6�MaM�h]��YJKh*QY�0C�r��&&�(��HBe�EP\����vQ�|�i���R=n�ʹ�7R6]��f�V�VjI[*I�гr5&I{�XVq�G�b�"U?�����.2&���#M�r�ݵ>�5!X�W��Ֆ@k'{�%���,�8)!�����]�`	{,�J@X���$�=�2p�o"���L�w\!���ٰV8m۷m��Z]x���wm�^����������>އ�Y}֮ء�;���wIȕmqn�q	m�^q{�Yw/P�����L}̶mLyn�������/�,�R^po�*���V�4ҊI{�S����=YU�}Gz������*XH'�
�Ⱥʁ\��K7D�p]cBzB�C����{�ֲ��:wL�m���m~������}�Oڗ��u_Ӈ0�*��C](�Yye�^NC�k����D
��3}�Z'�	�%.�jl��.����m1�=RL��X-�_���ĥ̥|�(�^~Y7�l�u��9�����,ģ�����.���Χ�+_��eSYvC~����_�%P�w��z���ݻ��x�⩤`$LV�����`��#�6�U_�]�DJMj4�6�xI�k�	s�3�S���F��i�ۼ�.J��o��x���a�����Hf�}>�ʷ�L�1��޴���>`U
n�?/O����d���p�*�r��r[���6�uM��^�l��>�s�6#�&��Y�/e������N3s�2?o�Ҋ/cBW}5��5lfv��ei/--�N
�Υ|+�	���%;}�� ��$E�j�Ν9a����U7\�=��2�r��eeӕ�㾻�捛��v�}����%�V�sp�=)�Jds*�����U?A�ʌ���|`@�����n/FEa���%�-�X�j3�^���12�����R���ת�N�b�g��L3Ym�:�Y�����tX�ໝ�7�(���c��$	ǆ�DzY�uudC�ےU�.*L�g�0G�@���>�/b��\5\�jUeB-���d�>��W��3^e���"�!_��kj�<Yh|����� �5I��kb����0U��4����!��#X��D����֧'��5B���K3�	v�n�^J�[�,t��M�a���� �qÜ�&9d�*��X�a&^]qU�H����R��FBNQ]�'-��"�Yt�V;h� ��B��t�����4\ץ}�@�+!��i�^�V���� TW��½��m����P�+�Tܼq�n��f����ψ��W��0A�`��&�خ&�C��	�(�.Apg��,aR�z�]v��)_f�UXWAPN�?��w���T��ӹ�p9��� �8�8�,8��Ŝ����ٜML�)��*��ٳ�W^��tQLC���L;s�oc����קh�-�t�"�-8k3X����x}\�V�j3JۦC�a|@��X��xXR���Y1Y� Y�,��p���LI+�j~zH[B��,�g��f���2�vHL���3��/��N_�Ҵ���ҝ�d����u�]8wZ� �+��*��Жr��
��*���w���yw-��F</�6j����:}V/�pך�_���k����R�617f�䠔�۰�m�{�ץ"������Ԣ-,�]O�֛�PȠl'mfaՎ�Z���m��>L�-10n��֌��Y�.�I`-�Jp�Ol<&���fo�U�);zn����ؔ����0i���.��`Y�Ff�6n�g�v
P����$��Xc�k��he�:��U�Ɋ�� '-���jMB�=zԷz�$�Ņ�!��¤��KX�M	&�����>�Li|I��+�@ed����6*�ex@|�j�����i�*�K�z���'�8�h�2}��X��N�YB�����~�8=�B1m�C",�8CV���#��f�TJz�D�<��|궾�i˜wSU��� Y���>;(3>��:(ϙ�4�pO�u9�6袐��"�O��L����<�
��,��X�W�:�"�B����c^�z��;��a��pP���g�s�3k5\Z�ʤD��;w�)�&)����N0V�W� R���KI3!�8��ӹE�����|,�`5�e�L���T�����#�yR}�RҤD�>	P�����6��	�1<ܩؑ�������@"}su��B�q�8a��[� �ѳ	�7o��MYK�bz�믩��)�bt鞶͝;�O�9Zk�I�m��ܸo�}���V(f%%"&FH��B�PnH,)w���x%P�A�?
��:JQ�]��e�x
������K/���XvP�w�%��PZ�L�]]�n�.Ⱥi�|x�{EW�#6AfyL��2h��)�(8��3v�o��������u	=ͻ�f!���.m�����a
-��++j�1%����'$�/���YG�fR��ll����nfo�^W���=�����ܽ��'8�N����/^�]Q�7l���&-��*�����c'mb�f�[\�)Yk�7b��;�f�ҟ9fr�U�,��^x��f���7��=`c��F��kgV��_zQBmXɤ��Ҍ�؆s�d���^}�a�=x��I	��� �>fN����r�����4�/|�i���3����מ|͞y�=��Y{��3��_z���s_�O�q��^���;iϿv޾��I��S��?��?���}�����=c_�%;sqI�^��|�E�����}Uy|���ǟ�^;j/yÞ|�e���}����/~͞y�E;~��ǌ�B�,m���g����]�tAX��!L�	333V�dCC
+^ ���N��u�B�&��g쌄KXT�څ����	vc�Ãy=Gi/뻖��S��|��{w�ԥ�=�Ks���J��@��m�Mr����_�$k��
M{�3vz�h���otq����
��h�I�9Pa_�@B=� X(��4��.%���,�x\��J2~�{i�B��u�����ɇ����|9�֟9��x�v�)�@��U���`M�,����,/��H�T��Q���a�:fs�Z�����,�A�!/i0�r�Jׯ2�U������T҆d�	6Bs�9ձOp"�+U�AYÔ)���Wǥ���>�+%��U'f$�ҦҺfTuR0N{l�^u�)�5ņśuK
�R��H����<S�T�dY�;���U��4h���+�z� ��O_vVAF	z\}�-��,�<�}�w��z.��zK�>	H�\k[_b�������3�ŜVŬ�lώm�<7mS��Y���-�W��פ �w��v�݇��[Z*���,��� �
s�B�ԬP/ͅ�ڂ�����bTDQ�Sܑ<&�$k���|ݞz�)wc2����|t�5Q=�B�[E�w����p�ƞN��D�����쬻/a#Xy�/t-{i�gnڸɅ"�)�$�r͏��2�V9zU������s�Ӈ:��"���+܏���h�͢�K(�+��?YC1	�Z�d۶��c�>`	��ԋeg�^#��[uh�#C�ʦ���}s�dFݤ����&�5;~n�JBc�wXM�����=7���\�W�,�|�]w���`�b�ڪ]�]�;�o�響0-�2ie�=��m@<�6b�}Q�O�d~����Z�	y96���&�.!�H*&��2c��,Ř~�������y�>۵u�TEYw_�Ʒ�3_|��M�,ݗO\�W�M�G�ر�3va�(>�P���|�p~��{�䔝�0o�z^k������5{���zw�N��$��*�+�Œ�;z���;v�����-*6��Q�v��		��%�v�͇}��+��b�κ���a���n�H�`"�0��en(��%��{Մ#�'�S>Ĉ�+sѷ��n�$ϋw*|c�c��⊕+�'iz��6���n8��Vʽ���Y;9�"�O��H����6��H�����$������N�$����6��R����a�{�����C��ɴS&�K�Q�,�t�13	5��4Y�6:u	��P�,���e�J��h$$�V�W��y�m`��dx2�*���oU!<{�� Si	`e��F�j��sV�FR_\��K�V�4��l����)��8m]���6������̬U/�Xu�5.�)귞��g��ή/,z��/X�(󽾨���4�������ݜ�7�6f.YG�*;��nU4ֳgU���V:�JΩn�ýb����VΝT�7�|��UΆX<�N_��So؊��z�:/Hs[�[c��*b2��4�H�	�|�
�m&�,M�N���n ?�"�s8��Ս~d�}6V�;menٞz��-%�%�o�l�&/�=)�T���19,r	���<���V�	�/�b���v�w*��5�KNT?���Qh�`�>m�+� q�V��r@�#�:��Ͽ`��$`��ڵ�w���U��j/S��^���Y&ԑ��:�.��}xOz~�0r�{�� DC�]0Th�v�!���\pŀi�CҒ7LNJ�$]��F��tj@9@�����B�C��Xs��Q����;��@��U�80StA�_~�ؕ�a�A��,o@��F��eT/	K)_����'��Z���������7���?�=�«���Wd=s���Q۶�&?���<2Y[���_{�d�����qϝv������.,�k�Oعs�����:}�^P�u�	f�}�&{��l�/��`X��s���OZ�w�:	N;OI�`���S)��+���+@R����㵪u}��r�Aۻu�g��
X�9k'OMK(�KC��?�Uԓ��8(�=�'��������쐥���@����
�9�+<���Tn��G,78*�w���$Õ�,S��N�%�d�����B����� ����{��ma��Zp��'�(��r8n)��}�Rҵ�<�����'�'��n�S%^��܄�>�G��;�!>ayB��d$��cބ҈~o��Nۻ����=��;vn^�q�29bܺ�F2x��;��I\,��������eF-'�wq�c4��H�?���ǥC'���G��l����(`4UQ ��>u�\����F}An]���n�u��\��%!�.7_��zxp�t��s<P]�V�R�ǪM& $1V�4Ye�̔�{�U+��`���%	��|��y[��Y�0!���\��."�ti�
8+&+0�gN��i�383���i��sEO�ޯ�;��'m��q[>uܖ�8j�u��H^J� Kf^�V�omVW̾|I�yZ��y��>s�U/=k	��fg�='��؞�$�J��g�[��ik,-Xua^m�`��%w�m3)���
abG���Le2��n ���h����v�;B���� �pkҿ1!j_�d����/�f�<q�ǂ�C�u�;}L�p�2	թW
S���##y����.���@���H���Y #��@ 7y�%DH�F�,Eg�z�WW%G��Ѹ�ߓ�?�*�^۱c����kn-B#N�����v�2�ǺFe��]��._a
\=z~g�;�E �N��8LC�	�V�n0|�u���w͕X�O�Qj�|(�Ji�w�@y��%�eI��>���a	��#P��1�^��מ�JYJ0�YK�lr4g��s��-��U�/~����Ge��8c[.WD�1Ѹ��*�_�B�uI�MI�*�6�ܴ�j�b�1�.Ԭ��E��+6��Ԭ������Y{���l~�`�ʪ,����2Ȍ�bEB&�pb����=,A��,8
�G����ϼ&Eq��;\��I�w���kV�n0f��tՍ�5��&�U[���E?��#�}�vmf�I�ꪽ��벶��_s��x�P�ڢK�0ڸx��\7�%U�7#�2ƶ�L&�%dd󪏰Θ1�'�R)ڊ�R,Hё2"��'R�Z�SBN�K,�&<�f�d7�
}�����m�?�m[���P��K�m��fr��z?(E���7@�T���dI�I����0LÄ�5�"vƣ�P$�H� _8)�y�k���7�w&gw�{�m޾��V����33Ek	bF��;v�hZ|a��&ؖ
N�΅]A^�G GC@|4�t0����y��h������2+���Ě�9f�E�EY�_�@\'WsM��Y�,��lV��Y)YoUZ{[�("�ݗm�--��4˖a[�Ʋ�Xo�r��u
�k��F�!�5K�W���¼�s���uF���oe�rB�\�eu͖��)�s�9�։���`��%K�/�ߔ��U��Ƃ�bSϻ1Ӥ~�_�~�h��v��T�˱Gu�z��,�6���,��ve��T1c��90�����10�+!�2O��]/�{Lφ~忐'�����X2�S=r��V.��"���GB����ZQ������t���s�O`�$���N�7f�@��U4�"
�G�n���OH��뗭pV�Ƣ�,*W%;�|�i+���O������!��Z��K�ԉ� �Te\��5A/n�z��UQeF�Q -���h�:�~C#�I�,��#u�a�掕�Ҙ���oNȵ��p���"�?�05σ�+nb���ߕ�;6�-�{� �%�Q��I�1��yr��?��*��u���c\�
+E�M�[�HzҲltM&Շl�7n��,�ѓ�Ɩ�g�$ ;#�bc��:`/��l_}��}��)��d�%�|�I�g�*��e��I������&P��Z.���pK������?%E��z�ύ�����r�0gצm�lJ����va�.��u{ٔ��H҆�ڪZ:.�׳q)���H�햒�q eCɎH�'[69�T�Sb�a(k���j���9�Ӑ�m��CFt���JE�1\�zW��l�]Ǩ�=5kvdE�A��ъ�P�^u`
\P��'�~�c�7!Zv@��w����E�!���^ɜ�,ɬ�6)<kV���#�;%�0���g�.3��<x�<a:V��vV!>�J(H]�+�rۦ�.�&�I�xaH����9s@tA'��|���~��,B�`$,�]ʪR� ��>�K;��!��(�ψ�.y\��{�DUΉR@�١d�e�����9b�J@Ĕ8�&+D�c�J��w2+��J7�J[Nɉ�O�� sk�iLL�;6(v1,BQ�\��S�{�6�+�5��[�U�4^R0N�����u��w6�a7-�n�^BY1�)fD�3�xvuL�"F��ʧ�Z;bG�$���^�XN��,�t)�/��]9	p��y� "<1����嬔��R�u������tY���2�^U}��Haq���1<fh��c��>	;�H1\��wq�����ҋ�aR�0�,�T$@��x'|�p����=��s�e���:dP>�}���N�`�o'H�o��i��5�-�OOݸ<=ϻt�>Dm�6��i�w��_���%T~�,�F�-k�W]�X(����J5
d�?����>�M��I�m޲��B](S���⃢
c516���`Rnⱌ������d�C�q$��SBt=,��-䬱����#H�_��p�es㲜��<�}�fESY��ud��r�I_`�P7,���a	8��XC1�oܶn�6KJ �JhqrLZx�T�s��M��(]Ru]�Ri����D?1d	��z?����9u�=�go[w��lLe���\[� ��H��^\3�@�P�	�1A��=(���Me���R~X��f��86�t6>6(2m�5Y���/E0*|��0f*C|�*����#}���HΚ����`2a#CC6:8l�ã���Z�쓊�~����^�҉;���=���<zA80�-�����J�"� �|�A������o&�."!��͙�a�Ƹ
3�0I�)��{�f�F�<Q����ӎ�pm  7�;�2���Ps�ffl~��ܰ>f1�y6���zi�A�����YOuDDz�QiH��#���+����1!S�y�6��ш$�آMZ�Ǆ���^�q,\����<2�$dR>�}⮊j|;��Ǆ�\�(pM�m�SyQ�c�+�=���=
�?\X������]�}���lE��,��rg۶osbf|`p�O�U�Ra���X���r��ַ�g��)�W��˯T�nq�+%o��J�X�I�|Cp���N�w��E�O���&�ti�S���]��d�ea2Naw$Q��m<���'j;�1��W_���x䷮�����@[��]�J��C���!|K?�^V���Ն��x��9;w�+�(��4�U��r�xQ�.��C�ז�o�iE,�0�&<g��z�i�w�t˥�`+*i�R~P�Y̏�B�0�ݻ�X>?�K�d��1��bԂ��ōu�k�B3��	:M�Xe�_�����Eؗ��������"'Q$܍IDL�b����|����Ҿl�]�ԏ�lO�֖���^2*kJ=��S��	/g"��Z�FǷؾ7�;�K�sLlɭ�3={���r��]�V��l�P��"nݎ5d��[,�%B9:H��R9�<����J�]�,AMQ8�?w�+�aʛwa#�୛���׷�cV��DC�e���;Y��U�v<v�U��uZ���~�&'�'~���~���~��t�1��?�3��?�c���q�я����]�{�[���;¹�ާ�'�=W�`��<�O:]f�Y�)�bi#b�7aG���*� 0��S�(�����fr���d��[	�a�iN(��3lѣ-Qd�Z�A��]�>ԅ��.�ab^g�z�]�e2˒c����FC�"M���*�]6�q\<Sc0eA�/J��X3�����J˪K@W�J�uJ&�J�u���:)"؈�Fz���rCY�أ஋���c�.G����Q�du�I���tō$�K��H�<C�q�)���Ń�= 4bz�D.�F�+}��
��v�*F���jJ���T��3;e���:���=�]�00���4Ah)v�_)�&��e;n�9���o4i�ѽQU�T�?��̙��$��.#Z���O(7�7
,������5Wn���]��D�~�6��n�#@C�p�Bh��w�����OW�X)�������1*�Ĵ{Z�)�������k�Q瑟�C10����dA2���z��v�qM0�?��T��x�,1���D��>+�\�'����t_��&�T,�I�V]�;Y����(5í�oa�b��⊟cW/ČC^u�Zm�Y�u�������	nMH�PjZa��T,�t)�kva� a k#��u�2�����d|�݅KKV@��$le�����|:����墭k�H�}	CJ�kq+6֬�굙bզ���u��Ip�dG��Iي����r�ǖj=Vmfq	~Y=���Z+[E����l2 ڋ	)��8V��T?b�$]��zVX*�jU�I�s��#d7 x�w�,�@�ff�Kʼ�6*��C�l�hg���;m󆍶��۶����v����[~Ķl�2���+�^��Q�&(�$���.K]x	��w\z�2���Ri&���A~���G��q`�8����ևg���k�zA��X��!���a��^��;*�5���k _OO��ؑ`a��˂E����Ϊ���b#�9AY�Q� �֕��hl�u�:��p9�����Ye{�����sI��"g۵[�(�5y�^f>"L��٫��J�:깮t:M�wc�J3"��?��WGe�h�����t+&����5�� s��4�jϛ1���F������ Yn҄��TJr3�(u[�xB̄]U��qi'^�U��շZ�c� oٝ�ό#w��e ��[��?�E'H���8q:ՇZB,Q���nMYC�w��!��� �$��[�nJf����H譋����
~]=	׫�����TM�a	6�~�����+Gm�"E��:��{a�>�β���
<�(,W,��ʣ�+�Aٕ�� fMY�E�)�ŒPY�`���8���+.Z�8e���;%Y%���E7��ʖ�խ�a�ւ��,߻`C�E[+�a��i[+����E��E��ZO}�z�Ko���b�UE1L\��,p���H۶͛�/�8��R��(�\�E�g�e$��%��h�	�����F,�7b���MB�R�@�]��ֶ����z~v^W�S�=[��s,(�Yo&o-��5�?+��}g�%I�ł��>��ǭohRe�yp��TK)1N������R��RQB�-ۢ�#k	�b)	5�\��)��&v�Ǳ޴��m/���q���%���C߂ѥ�O\�]��|�lb���m�k�.����m��d�V+-��@Ɔ�8ȸ�6m��;7{9���AH��w�I�1.��$�BAuQ{�4��G�_�[�k�RC�|ጝ��l�c�-ٟ���bz$%k1�p��F�ӟy���$G�P+��3~9��$��Y�U�70(dG�Z�-�6�M7�Q1��g"�����E}�է>J�,�o������b�eO'}���p����.M�h��\8��O��hsd:�B\ʁ�/�{� ��������6gDݫР��4�9����/��E�����֓n:o�ޫ�zN����E'�1T'���a�G�6D`����]�Q���o��k�Y���|Ϫ>�d�';�pb�Rɋ@���� A�ߌ	�G������ε�ܲ\2e/�x�^��'�o�M�{�*�� j�«>��RY���E���u�	�5�)�!ħ�>�ޟu�9��QR�<ǅH*~���K2h�-��$�z��_�ǿ��뵽{�(�rށ0z�d�3����n�PWڭ;@�y��+ѕ��Ú���9��Qh;���;�8��!{�L��-�Qٜ�}��E���÷��l_~��B��1F`���hꂰv�.�!����CE�LQl��:����N���7n������#?�A�`��f��y��{��[��������G?`|�c�#y�}��o��������G?l?�C���w����;��>��}�����[v�c��w<p��}�������w>x������v{�Cw��>�^��������؇��{�#���;t`�MN��2-d�0ľ��c�ԳG-����I󲯲Y)i-	8�!��Ә��l�;�Ո灍���<{��o�`7߸˕�7޸h�����O����zoN�L\x*���KAn1wB�X"�I��_�	Z�-�-�TZ���eY<"&���ǥ�#����R�ɚe�DV�	]�9��Z)�}C�]8c7ܸ�F�F��g�m3�i)�L^�XVV*���9Jz�v�����m��"�d|������R�E�>�zt(cy=����=C9���#G���+n]�"�l�8Cc�?[>����TyE	��n��6l�"���^�hgf9�.�w�{�.��^�0��B6�-�n�!�~tl��]��B�Ұo����޻I	�B���ʃO8R��Z�ӫ#	N6Wg��];�4^�"�:�+3P}|w�^t�б�?l���viҾxKww�؅J� eq�y\i�y�9c�Mz"���vd�L�Ih� ��ϸ$�Eʕ_� ��:��λ��H�w��Ƚ./6l%�CL�r;Ҙue�1��
n��2[���4�_Bl�*���2j3{h2�:AT�K� ��|Ӡ��Ł(D�M	��w�QA(�2�>�244,�N�[�3L�V");��w����l��MҬUO�E�X�m�>�$
���eO'����UŽ-�y7�6箑^[X��n�l�>22"�3C�(=�x�=g4p�0��6�pD�6z�<#��^!���HP~���"t�&Չ��ʕ�-dK3����yq�ԃb�t��i�DJ-u�ܚǛnD��O�7�sjwV\h�������lH�V���B�>YX�CvϽ����}���{��n9����fwܼ�����C~��}�>ۻu�n?���9��n���r��v�޶�~����s�ާ�C{&�=���n����c�Q{�v��=v��v�-��{�;��~�L��`c�����¿ĪZT���Y.���!�����RK�&E�0�,U8f�%�ZR��<��0�8�F��616��Z� ��J��If𠰁��,�T��H��mK��D�-	�؃w�`��>f������W�}ۑҡ>�o�b����N�d��.Z�v���F�WC��=:���Q����yii��D�`���,�$GZŝ�|b���τ%H�IaawƂ�>�N�#ePW�A�R�������ST����J����G����!����4։_f��ʳ~�@ࡡ!U6*������31�����@@�oYx�|��Ǆu����*K����\������YP�I���啢:W�@h��K@���gkk�i��y�}���"�!.a��q?���'�݈���Sk}@�����5��.��h��r���'��hC{[�ޞ��՛v	�>�b[�[��n�%}!����r��B�����!�I?|_ �N `O�G�kA�(B(E-������Nrֵ�FL��!k6�K����g�/�fZ��eJ��� Fp
A��	��Hy|���߁�0p���؟���y�a	<h�6]�S�)G�h���k�Xy��d�=Q靫�+y��+��_��fU!�1�}�v����W_}���3;����K
�C�5�uY�	�0ڥZ�o�B�xޭ9���ӗ���X�?�)��4��2Y6f�F�z��y}�P�R��S�7�GC����!d��!�F��U�CذK�OC_��{����YZEw��$1͕I�X�{[�%���������+,OK(ͩ5}�0��8�ߚE[-�*�Ek���A���8.(߯v����)	���sX-���-�7�Z�zi�Z,N��M�ۖS=R�Q�r�����.�S����Vq�)�)�j��>�������?lo��v��c#���'-��Kk����Sµ4�T@A�"@c���{v��M�.�Ë���?�����GQlH��Ž6>>&�e�Qش�?���iT붸�b�Μ�����[�&�1u����a�>���W�F�צG|#��,Cb#8�@�Mߓֿ����H4n���8�i�yc` ��Pp�������#zx�M�F�︜:%7�u�o���+TK�xm �o«+	�-
Q9�����UV,+���XΆ��if�"XZ"�&�7aE��]��[Cyy��M+f�����`RT~�c���mL�㊺6�;���Fi��~GiC�ʇr���Vd��F��x}]Z�ƶ��)����P���BG����&���W�JpA�~��H!2�&&�E��Byb>� .aa@h!\$�����#��b��l��)D��#6���#BE��a��etBfK.4T&����J�L��7P�}"!zѳ+����j�\Ϸ� K�F}���R���������n����,�1p����m�s�Du���z��^�OJ쏱T��^��i�T�����9;z⼘_G�;��p�ZY̱T��-(����il��D���e[*��o�(��>Eq(����_�B�� �©	,���,^��%e�=1s������U��'ldLƄ�K�֗����BHp6o�����$���L�~	5�_�V��ʼ�KV\�5W��211lY4�A�4u&�5KRH%�e�EJ�ʖ�T�fMJv���ͥ��RT�K�q(e��XG�z��Q�2��)�$C��>sqPےꔬ���OEX�<�{J϶l�h�YkI����e�Ǖ�@O�,���{]����,��v��}��m�KfrJ�:��+Q�ɕ���x���(�`,1�r"�J��Z���O�!�a#����|vr�וK�'В�14S�!B��K�� $�#��.;�bX� ��Y��ѕAq�^������>f���?�A���bRI&T����K�����L���R$f�~_�A�YU���|M�;�.��Uh]L�.f	��ҖL"�ĲCţ���J�ߖy[N�m%���d��"1�g�̀�y+�h
JWH�bi}LD1��>�ZzЪ��!��ĠUbVV�ĸW�X5��ǐ���.֧g}V�EWIH8&��&ZG��&8��]m!�/@���0��J �Q^�+��ō�����P��F�����4���$� ,�ٌox��4KI���I0���!�Tt�,�`��uuhy<W�� �����op뱈�i� �&�G�!�\��Q��Ӡ<^[|�-���|N�}�#�K��3~"�Y8�Q��3_k؍�P����r����a��6�(_m^��ؘy��ݶg�n)5K��;s~�~���=�����=��I{��{�ܔ�T�/'<M��r��^�d�g�lzaŪ1o�Pfx��;�P��_�g�N�ѩ���d9�����T����O/��K%�[Y��N�bɼ��~W-i��;rz�^81c��_���U{��JX��k�e�o|�[��h{e��l�_�K���J�����zr���Վ��$L.���,��!���Q�}%#3�*�K�`J�0��Xk���d�
ΈrJ���I�&d�e�o�R�iߟ!Ƣ�o?��=��׭�U�e��%(��=,>آ�N�n	"�Wy�)�#�{(߯�G����m��(���0D �9t��u_e @�r9��*���K�v���/��r�.3k28Xz�b���l�P�sG{T&��@�D�߃�Dv���b� ��Ë�o D.�(PÞ�镵�,�3�u����}���7���7M��/>�F��|����!b(�F �C���9*f cJB %B�8��a�h�������g�*�����YISR>��֫<��<�>ęu��We�V$��g�/�m���7���
�W���Ksї��Hc�4`��������<j�1I_N� b���@!�L.|��O����l�C`�T� �~	�Bѯ��7���T�O(�v���;	m�N�è�}Yݶ�Fvn�y2U!�3Bqi�M�˂�7Ւ��d�9���̘0���W7���7U�L���/k���.aR�nm��Rk��FM2�~����6n��&��>��X}e� ζp��a�6ؿ�矰͛��o5�B�"�?�x��a\P��逍k�C���`�̰�ҹ���M���r���O�s�>��k���ުt���l�p�ތ<	�!"�HX�/����N���gDW�TYꆗ�<q)�6U䫴�AN�|�3�w�_��B+�`��%-;0l[v�#�O��?���i�6��G���U'⺧mL(��n��׮p��+�I�wiqXf
s|'�/���_�'�ē/ZvhX"B��J}�d^�=;7�捓6:$fY)�Z�'ψda��m����m�v۸e���0k��^����Xnض��a��t@�T�
��+Țصm����������=§���vqnƎ�:kGN�76�߰��&6�P���<��K_��=���}�ˍ['7f=�!۴e�q��k�|�zYJUkK�ݵߏ9J��[6o��s'���gm�`�~�?�C�+k�m�f�:~����?���Ꞽ`Ա�ɍ֛�Y�������9�F���0ٲs�--�Z�<c?�{��G$�j��7������-�S����-\���yY�U+�.����w�J�cu	�����jI�)ؠ$�/���n?�#��y������k�[^}�'o}��w~�+��c�6���{���,<n��7�ly	���Y�)[�U|<oۖ-�q||�
_}�U�������K%[ZfhQ���J�����X����q_��џ�I��̴��__���|Q�q�m�'��}v�&�_a��VU�Z����O��_���mmlø=�ҳ.=�-'���9��b&jT?<���xv����.�L�	��'��Y~��>��A�U�Idx�SR���	����ڰ�BI��� ��cY�NK�V��2����E垵R9�щ�n}0�)b��f��ۑ4
�ܻ������5p�¯}����q�(x=����|��0H�3��D[n��:B�9!�~�/���듖���rӚU1Je��!���Z���.T�?�mW,Q+�c��[N�_��߲�[o��{��W^O�,�e;��ڿ����M
O�1z	��! ���s�xM���Hh dZ�!��r����������K��y�!�H	��#��x�)�{x���Z���m�G\�HP���޳bIYF����o����	�7������V�J([�!�"��5���[;]��C�=s1ϐ2���^<�T�x�M�?�G����ӟ���V^��0�h�������m��a����?��$挋.&e7��z;f��wټpv��nI�j��_u6)|=�X����x�fΟ��zZ8��2})���ĥtw��I�|��2鸍�g�_ڱ�^}�t^B�or~EZDp�����b �,�o�d	.��KP�̞���c6�����O�=�6�a�v�R�~�Sj��ʷ���mON������j,������Q�e���VY�U_��M������}�}�/��Ǭ�Y�Z�j���=��V��c��%�	�H��_������-K��^,.�5�T��տ�3���՟��G�ڿ��ߴW^͆��ܽ�2 �����z��t�7l��x�:ʳX,�D���aw��5Y�ꑑu���[6ۅ�S�ۿ�)��}R��R*��xW%�7I>�Esj�Z�^�ёR�c�韵�{��M�����}��~4��|\�v�F��b��g1��9����(bC�fSX����ү`���~��B�V��������������(�'��?����,�줥(�$b�{i)�vC�W� �K�6D荌bN����5=+K�+%�	+v���1nK��% W���(
�
���1�7۶�N���uN{��E��ps"�z�fkW�i`E�3b��+-�L�K�^ԻsҜ�*^�6삐d��j��m[Z�V���͵/-U�!M �!6�|X��z�;�u��C��B""km�~���Ȃ�P���#���G?��)�]��� ��th]q�����(�I�|m ?��t}'!�1Ͼ#(͛��:��+|��fa�������`ǆ�xF�Պ`��Y\�K��A0�����	ј���>D�b�'��N��&e2�6(!�Ɵ2I�	d!�ټm��Mn���~Z�Ħʜ�T��a[��x�*+�z-=���7�`��FYiC֎o�xn�e�n��7ن��Zvt��'�YnL��M60����~	�=�a���������l���-�26��Zbl�I�Y';f�Ā�%����
)�JQV]O��`00!+m@�Vo�
~��&\���И��v��9+���R�lG��R��g��dD��z��(�����v�X�?n��m�}{7�*ﳷ<r�=��{�"^)���쬄`�6J��ڲ��l�d��};���耰@})�g�G/�œ8%˿W�9���3�����3R�g]�|s�� ]��Y��甜�g�ؑc'dH�j�z����⋯�fo�=cO�j���~Ξy��֛>k�/�Τ<�����B����6N��7����C/�~>�b?5,3�Fi��\�vc�-�!�
��0~r�n�A���+�+a<�J�w�K� "������p=��E�f����=�>Q -���(m� ,*���+5[P�+�m�԰iŋ�U�(�fZ��I�%�&�-�w�*�#�=�.U]YXW�|>��C����+3BeK�]L�J�'�-{S���n}䛖���Q&$�W����Y�+��?	�6WE�eu|Y�_��~���\��XD�Y���=
�;����د�!��(8���U�6f����aQ���Btl�-z��E�b�Wp8�(��}��ׇ(=�:!�R�欛^��X�BA!@>��J�>wܪ�O�����>
��0	&*��D	���������ō�����(�CI����9����2,x"߬��w���\�-"+xT�fޫ��	nq�������vv�b+��U�=V���rAu������^65h��1�Ϡ�I�,13�]ǭ�JYe5a)�����BŦ�����-T��(Z�Y��XXK8�]��dV
q�,����I���mz�nK^���q&o�T�X8�VDy�Kr�;�ms�N<+A������q�(����lߐ��S�mvn���3�M�����X?{��z:�~�զ�/�Z�?f�z�����g����a�������/����_�{���lVeݕ}\���>��������_����O~�~�?n��}�O�5�#���A`όqb�xR�_]�8sP/i�1kql�yU@H᩸p႔��UU��������v��	;y�����k�����}����'�e/���/�b_��Wmzvޏ����p~!�h��>$-�
M���q;p�RY�9	{x	x�@e�2����e|M���4$�bE,:C6��ېe���3�&���=�~��s��P�笑�}҅o�o�נ���׽�*D�`P�2�ߗ ஐ5��!�!����%�mM�#v�BhY,��Ȋ�)���I���P'��z�&M���"mnH{n��i�_ 3U�ab�����G�G�g�"� ��z��#�l��T}G�Y'E���W��H��w�H�*-3�?�ۀ��>��	#�~���H���E�zI�#��t�14��[R>���Nļ�6Xq�>�F|}��k�IIH�,��)(�n�냾Q:\���u��xA"�
e2�iH{�����vd���/�Z$�"��^L!��B�P�����W�����	��p��7uf\y��͖��QKP8��n�~C�t�Y�5��łM	� [X�鮉�D��*1���ID��"R�Ѵ,��u�p�Ya�0�t|���UZe�7�t�z��?	�ތ,�L����60����,�L[���Ov[���Q_t���JPg�{�tƧǧ��P;�-���^�����u���	YRF٣��6��#��]��ח�u�,�����	��k|9�A��{������1a�|�]�������cS�+q�[k�P�l:}�v�ضͶ��T�{[6�K�"��7��I(l��)������� �eW��o��F�'���h(��h'
��ܻ"��t���ϻe�O��X����������(p�<K����6u�+e�C��|��'�/o�_)��>�,�'�� S��ݪ��Đ�#�$q�g���,
���/���x�&&7��Z?|����cb�k�6n�`����*	���l�R�7or�D�0�)�;bĪ�
W����Tj���v)���Bv!B�#�̊�"�=�[	}̑�(Le��i��;2K0���Z���x��&e�QN��� ?���,��;֗��L�F��^I��)ț��&�V��\�6璶�?�A1������(ڌbCH�1:>a�VVd;���%�1 ı� ����}�Z҄[��5e���'��-�3Y2L�QV��cs!�+
��	���5U�'��Cx�[%���B9! `��6)��|�&��J�.�� W�-�j�DX�S�5��s,����� ��^�T,�hM��N>�}�L�V�����hJ�d���<;	 �;�ƙٟ��5ju۴qchF��A�0<
��Z��0���2
K�R?��)2p�z
]%VU,$��g}@�_�	�W�������%�f�q1H�]�ۀ���a��N@t��es�t�[��O�9�%[и�)py[�,0���"�\��;����\(�W���#�'���8�F��frFCBݪ-)���Ukzl�o�6�6�6�կ�4��64��-)�l�E�H`����� {��E����=vX��\`�LC
�ZaZ��\�hT���)[�;c����D�-�gU�;f�cyk�f��2e���[��T��n,�V����U���Y���}��,���m��e�6۰Ь�x�V�ZOe֒�>͚%�,��e��ŏ�K6>�P����U�3.��_Bp���E����l�ײ兪]�^��.6>�Js��(P1`�R�lV����������e��29'O8 zp�~�,��E"��#7�W��Ȓ�R)���ի6�0�zL�z\P����ڶ��lo�=%�y����������4J���z�G��I�O���,�;�d�g�� �J0�F�����Lb#!(���L*�
���� �mhAD�a8Q~�<�E� �*���u�2ڪD�O�����n���ȊW�S1z�����E�!@�1C�BiH������T�=�T'eP�����n�R�զ�t���8�E!��%k�;a�SG���s���3K�>kE�ʉ�l��u����Vta��/e�b��eNZdV�	��)͓��A �W#4&��)`&&)�)����O������C��X����5��B,<vhp�/a��T����
!zr����['�M�Lu�P�hp$v�XB�$!}�����g,��=Q�X��c���kN?w���G��4ݨd`�5�y&uAx-0v�l�05u�w�A	j��c�@p��e�>
n�)���P�h��}�Y��ϯ�S�ݿ��n��M�:�7!W���M�\EѠL�_�A�(�1�vU`	��	x��>�ם�I�pQz�_Ѹ<�]M���M��>G�������Ĩm߾]Ve�A��[E�3D<!LلѢ�r*ދ��F�������Za+A�N�7%�$(���j��� T����#�u���L%��+���)���-��61��xKB��d�Ғed�F��*�m�6����f���,Q_�����:U�P22Ы��o�l�D۶��[N]9��)�Y�Y��D���H>񖆧����l�v��b�²}��O��R�Ku{����_{�^;qFm��9�,�挾��'�����O뛧m��j�KU	=�W���Qi�b]�V��e-K&��d���`��ˉ71�� 1(2�-T��w����K�z�6dbΤg�"�g,��焇-�P��s�b(����.�D��"�t�������ietQ?&�����rO����[%���*�5�˱���8#��-6�D��x~����0*H������+h�!?V�6ZQ����&@X�/��
��w�li7�PvB���-*���˚��雽�A����3"�;&+q\�:P.Z�4�sO}�N�����?mg���v�O?eg?��v�K��ԗ��N}��Gv�`�?�v�Kd�/~��N�qY"�qi�����Ǧԫ"F�X�v��s}w��W��^���j�÷��~q)�����W�GA�^�,t��)�<�� ������}UE�~D��nf���b�u}�=����ؐ���ǈ1��\L�o����L�_|}���?�#-�z @w���|�Y���U8�7KEDKޑ r�T=��P���h��M�}\�o�G�2&:����:�m�e���:�p��~<Ip��tw�`���,W�}b��034m�������x�@�c���x'���|�g�^�.��au�IE6�犕d�+����]0mo��9E��I(���`�w@8���~�t��7�75��Z��G�X����k93�C�^Y$k�U�_��"B��헵��5��I�0�����>�Z,X�D<��-{�ȫ�pްR����F�2�d,)�I�:���O=sq�~�w��~���C���������k�/~��?��߷�_8�1T�&���W������>��f�����7����O������we]_%�3Y6��'�+G(��63;�4T~To�k��dM,��_�k��
�}��(pcv��Iۼe�MNL����m�ۜ�H�*8���
���)��ѕz�)6�T}6�&/�c��M`�v]q9%2������>kd��ُ-P�Ė�Vd
����2̈́��g���N�L�!$v��c�B 8^	���Ir�%n�)�������W�ݴo��P���=�֑�ޑ�%�\;̳�N6�&�e����E��2͛'��̓߰��C[������m��[ϩ,>s̒�G-5{Ē3G�����{�%[;�}��?a��f���6��?��o}Y�_���y�69(-/-s�%bv∠���	&ݍ ��5Qj,��� ��6K�����F9�}*"uH�e��PZ���7���_`����QV<�f�q!j�΋��"��0������DHA�0�rY�{W���H(;0�,1f�"��f��4�B/>���yе����2Y�:��ٮ={|�sRV�������I�"������������G�k�=p}���1����ҾI�n��9����*/IL���f��3a��ب�3�D��'N�M��J�[���;�F���m8;-D��"�Fz��3q���M�(�u��[��B��u�[i��3��d��Yc����%��=E��y�����x��c1xB
f/>,���{<Wm�'��b�e�N�zs�(߰�y ��u����	_e(]N��~��.���Z�%��t$��������*8��ʿ��u�]յ��=�>?�O�b���t~���s�Nٷ�9b��5����JӞ|���y_+Xj���SS���vVB�-����R�/�v��i��x��94�s�|���+��;o�}�:=�1����.���s��ŋva�ˉ��%��Jտ�@D�ǝ��bvZ��r���5bR�������3V
]z�R�PF�^VEJN�H�Pm2���p+Q�
Ƃk�)�>�r�&��V�x����BQ��"F(
��󽆐z}N�6O=���f�����E_�XZ�w(��L��j�zV����_�����36��|�Iˮ���ֲ���lc�a����l8V����"A�bC�˷m`u�zOY�ԋ���v򫟱�O|�_�Z��Z^�b�@��֭+��H�TWMu���� �.8��BW�\�?/Di���BQi�%�{����o��3��)�y��T��94N��
�����G�s`�r�����#lK�$���c� J�Bg�#V_��^+���Y]�l���e}
����� �#��
��&��o����ъY�R���\�Ip3�ٴ���MDH�� �op�u� Lq�-,,�a�(&>W@���sqtM�;�W���%��є�k)JA�R�֮��"���Z%����XsVV�Xb�&EV�L�c���}��B�����*�~L+�H�*JJ����lv���!���u\O(�);)x1�T�h�YC�(�1����ĕJ�V��q�T>}���s³d�v��k��aKf�x���{2VFвE�,˖�M��ue�����o�R%i�X���-7�̽��j���X�q	��a�I���q��Df�z�}��oaq��u/!�<]��/J0q���¢h���׌�E!��(���o,z�Ƭhxzz�Ο?o�3�.T��M��<\M?=��e�5�#��p�!��,6$w
��x�����4��$����ޑ�"q7�:
!�(2тASw��; �B�-�E �l��}�
Ȭ_�M�=DW�_��:�Lad�-��-5�KXxI��]ݔ�v��lȖ�&�R]��9*�x�@�6J�$.Z��Kv陯څ���f^��O>e���6��d�%˴-�Z�XsQ��koQ�T��X2&��+�,�S���-�^����Y[�=fs�~�.=�u���/�"<i}�%�eٗb{"Y|j�O'�pg�<��ׁ"��O�W��]��]��[L�u`]A��!��rf
|]�з�
&5�#_�QVH�rf����� <ǉ�!�7Z��D���uǈ����Ui�Ѿ\�3ۀ��spQ��qS��wl�)�dMBPZk��-Y �I�c-'�(p�EX�A	(�?�OW�a� �n ��+B�z7��o�&�g���WJs {�N��V_�ߎ'j��l�۶m��Ǣc|�$�}GW�m��;߸A��=��9K��&�E�6(D0���g^�u;��q	�������m�fk���C�5�\4�Ƶ%��)�"eӅZV���]��jQ�d%��.���:e�ڴ��-X�5�g�Ś�0Zbz�G+Z:�j��}_�5)�k�Y�:48�oe=�f�{�gO���1��z���d�%�:��,��\QV���,00����ē.�e��Ldl�ڰ�O_�3Y?�U�8�b������kkI���[:7d��ˑR&�i�f�R�1	7����J�NO/�R��͌���E	=�Xvh�5{��\��lBC���b�[Ʋ6�����P<��I���kՊ/+8s��]��d�zNg��N@��k�+^3�7b����2>>���>�'a�����}F�B�mGb�݀����z��/GPa���tZ�G Pb�Czx�c��w~��U�R���KU{�ش�oqB��	�5W�I�Q0��Ajk�h4{V���0H͚�[̒A�4�����%DO��M���pʧ�Ċ�Ph0��t�H���As�2wbj~���*�%i8hB����F��3�X�2�"C�5;�dW��O�lC���⑗�̷�j��}KB��,�.ZV���Ƙ��92����E�b�quJ�L!0;�����4���?����U�۲|��l��9�zY���&�s�`�ٮ�CQ��H{�lqm?8h���i�_��`�<hv�`G�zM�-(�%�p��ݤJ+���y���C�R�'����
�����r��`7���>{��c꧔Mn�`��P�?&&\L))�޺���l��	߇��X`0of^��_<��p�����{��1dU&�f�
~�ئz��ғO>�<��ܙ�ȉͫ*�.�bPZ=�����8����»�"����,�A
0��]:󼨮�?���ދQ;a8\]�V�NH�g߼띏���o��70����7톖ݫC^�@�[���n�!�\��J0
֤�h���e��ן��V��nT���m�Ġ,�]v��.۳{��d9J��I1�${�������mv����{�f۴a�޸���M����P�߸�n;��6��l(ݴl�j���8����G���[���n��[FEg�ϝ�m���iӰmސ��Nؾ]}���撄dQ��b��uX�7��S[��t�M�RQ�<k�\�RR�:�Y	,�~�m���ջt6.jA|"kw�u������Q�0]�V~9K���D�V��+�5KbVe}gR)�,SHۚ,A�,��<�o1�ib�ޥ����۱-�R�g�F|Z�5�>D�C��uxlL<)!x�sI۵s��z�&?���o�=t"�̇�T6.I����	�Z�(��W\�|ބ�(P�sǅ��E�(�b��PC(f�9�a6)B�����b�~�wwy�{��6SZ�5����=7�|\Jԯ��/}'���O/ګ'gl|�vg�s��@��h��� �a��O��S�!�\.������������G.<��o;d���F��������C����ȁ���$ZJ�T�*"��
�� �T���S��W��.�mS��[[u��j"�#�g����ߴ3�=i��Zo�$b��`JB��^E]c�6�q��#!a,�!�+W,ǈI)���ΗDftl��kyz�K��	(	���a4_ή*�?Xc����������_A�������'#QG��w\���#��AwȠ&$�����ߓҥ�n�O`�����9���u�x�2�f�kE;�o�:o�u�.!�5n�����4~6�e�q��h����yۍB|1 )j;�3X!f��Y��fe�y�ip��F�c��6�R����#"�����	+J8��$�urD���<��=�2�g��81��ԏ�O�W��צ�W���.�!_��Ee����+!����(k���J{��G���/�R�$�oR0R~��C����������'8})�L���`�.���g��|F��>�i�`_�~�G>d?�c?ho�A{����n�춃���������m��Cw��mv�݇=>x���7ٝ�%�n?`�w��{�.	�mv�-;�;�H����w�n�q��y����F����v�m�}�|�=�����n��>tXio�{n�ew������;�؃��<h����RU��#���A�eSR��D�M��QORt�Tj���8+�U/XN�ޣ�a��Z�"k+eG����^?-q�x��R��E�WiW���X�^0)T��1	\v�����Tb�vl��M���o�/�f.�+?�> I�Sd2K�P�(��+p��ҷ$8M{de�r�~��^[Y��W_~Y�f��!\�8��&)a��@�~� ��^`��%�=z�~(܊��O�o&�e���iVx(8�ª;0�؃I�m��5{��6���%[C�ݹ��	Ɖ�Q2���Mg�08e�qфg�zq���s�O�H`p�@%i4e�V�"#�j��3y%�=S�.��$�wD~9��	��Pg�yH�V���g뿯�W��^H�jC@{G�ֺp|��v��/[c긍d:6���L��i�'��&S�&'Ζ�=��Ҥ%8���?��u���&P�&��IY�� �Jc3�N�aI_��*!ZSe�`����y�����gl��m\�?��� ��#�|��.y�F�
�V_֭�ۺa��|�QB�����l���8�C�B���w��!H���!���	PZ�Eu�-J[d�m�:��Xs!�L/���Ҙ"xf�q�S��.�����q%����-�,wtO���;��2F��M�:��(z����q'}���Q���#���hDy#Լ�j�㧾��D��
]��^�k�rDs�T9LR�HK�Μ"M�o����އ	 �ؿ;c��x�r�p�~��u!0�+�>�v������v���fh0m�<t��u�>�"ƕ�7m(������������IVٰz�ƇR�J�66��|��D�6)�y������ݮ4�n���o��vo������6[�<;����`�r�5Y��gZ���{�v�d���7f�ݶ��{���y���<a�eY4�X ݶ�U�5f��y+�\���K֔ŇZ�2ʸ��p��wV�E�(�t�7���L���E��[已0'!X�5WV-�w�H�g��e+�,�>��FA�U��jњ.L����|�����g���o�׿�5�OtͬU�m)��}��i2e�-`80�MA�⛢��!&���c�0U���gZBs���]�v��V���s�D�F�]t%tH��2k:�IQ�<1�p��>]Yƨjׄj˸�|Ǘ��:���v���}QEB%\�UZ���Q�'�PR x��c����1$�遗O6�U��\^xqݠ��+o�J�� ���]/�Ђ���9*8'$�g��_��c/ZJ�5ї�!i����,!�=�N�\�5i��j9Ǉ���������Q�������n��{v���l����}����6:�g}�bU�l�"��r��GE�j��%ʗ���k6���m���֔ H�Y������Q��7�}ND�~��;�@��o�-��Q�69:*z���r3qE�@t܈̚䜬j��-b���C���`�a+�u�NļQư��U�s%r<8�BD�1���������=���>�l��%�ɹ��(�[��Q^���D`���u�6xz��]����Û��D�	!�*D�*��l_����|IZ���{�;n�|>)�!Bh��	�������H�]�2���P\n����B� �ګ�JV?������A)�i�Ӓ21З�v��U$�j�O�L��:��Wi�a��X��Z/�[�U�Y;����V�zE_���g�z7գo�%�O]yJ��o��T�V�|f�[�jZF����Hr�pއ�,	�v����2d9�U�f���,7�O�R�K�NJ��S[:zo�4���Ka..ͺ���ȶR]W�!wMmm�RBzVm�9���`ب��T�d\�P�l.aÜ�0�d�<�c�&�7��͛���R{��"@�KO֜�'�R����B�5r��!ۼi�� ��f�O���H�A����$@�ᄄq/��!��@߈T���c�נi�Cڨp7X��(�k�*�3���E��҂��2[.r_F���> s*�e ��4U�W�n&4m��lLiA�@~�{q���ӕ[ ����7Q |�r��.x����bj�p�����Y�>�(�>���Ā�h������׿l�=o!�PV#bkT+b 5Kd���<"��D��c��w�/����}�m֟�[eeIH\�lÆ۱c��ݳEBo�m�6�mӘm�1YlLFa��m;"J|��#�yoͲV��N�*���o~ɦ^y�"�>�-���>B���)�k�=����]��w��~S� {��6`�0�DD��Z�s�e�S0R�-�V���BZY,�/��8u�;~�*�%	&�,-/�*\/�2�h��$&��+0n�d��ƍ�C)��<g�i�_Y.ځ��]�.--�6S,Dg�&�2£%�AdL�O������=\��n N�3�����s=\	��u��\��S�%X��
�CU�K���$�v���b,Sܾ�����z�3���C7�0� �@����łE!�`���p)p�-9z\�[m�A8��Z�ˌq�>aM��K67=/�gYxP��l�^���r���"![����$�:���eն�`�t@�+V�ڭj�[S	ݥz�����rUV��� {ue���٬YZ�X�1�-�#�g�H�edE�����k�_�8JmBJ]y�/]�FA����^C�nƑ�Ѿ�P����X��5���$��Fr6�<2}�)�''xq�lK���7��m�mÖ�Rn���+(~�F�6�?��J�`Zu��[��*�0;}���P�(����82FX�%%�|_��
���J��������&''��ȀR��(�6WC��s�Ik^W$��둉lx)����ߴy���G�	8����Oƒi�����O�珜���I	����]R"I $_l)��:�
�w�z�\P��4GD��
Nfĵe=qD{q���5ˉ���F#�}֧���1Ht*K'`����Ų?��K�YU*��bM�7�k��l����4,G�{���+�zuRB�m^H�?kv��/۷?��Y���C�[ښF<Y�P��N`�M���@΍�9������n����f����>�'��o~�ꕦ�9�PK���k����k68��}|�� wl���'�2B(���d�KlF�����,���G,��k����I;mi��	���w�Ju�6GF(�20,��%3X����9��2ld������\�S��4�(�+/�'�PW&�@�Ҫ�YwÞ�x�=��׭�V��D�bʩt�N;im���7���~�-��w;!cY�-V61�<4K�����!450`��;�#�G��Ȫ�$.jL�bi������C��kG|��ˁ��TJlI�gR����4��!a�Ƽ�E| �R�x�y�b�^J���i�kˤ�_�~���[0'-�9ru�f/H�}Ut74��2�V�,̯83�؏���i��kkV*��3��[��Sά�q{W~U�G�W����\FP�Y�1��C%�9�_H�ķ^������b���G���R:ԧ�����>�;yr��ꫲl.����1{�g�ȫ���ًVZ���̢������7������}����7l���Ϭ��7.ڱWN*��M���7�������;��Y\,�fΧ�8g���+�`�ϕ��%`��ڙ��}�c��e"Ȑ���m>�fc��׭VZ������c�����c_���BQ����;o�1L��b�R���T�Ξ����e��!~ۗ��M���K@$e�qlVK}'hKX����xE�`��S�B�NL(�#cV)�ߚ�ĺ��j�A>�.��Ŧ���5�g��o����[�B���Y���e�J�R��'�xqZ�eYu�s7c���������P|8��]���q���N�4
o�!|;66,�ԛ��^IIf��>����ڎ����i+��>��9;7S��0�g���.�:����0����!D��D~C��A�C%�c)?R8���TW��B`Xuَksy��H�I����Ъ��	���W��CG����<	ܶi�bU�Y�4�Y�f�8,����/���c��X�\�%mDa@_��=�����T��HP�߽�n���q�)B4ܑBN�(m�Us�Z�eؐ6�V���6l�,��7no�+MmB�Cpb���`ȁ�X~0%b�Z���i;���v��,�Z��Z˅�|GLFW�u�5��Cgf�{�L?=�v�}�!�`]�������7
Q`�M!/cE�"S�`ԒBմ\~Dq��28�d'�GQڮ�x�}���+u�����K|Xbh�a�	�PvZ��84Lf¶\#ݺm��ݻW饅J�Z^.�h�1}��
0��@I��J�"-!��*a�W}�.�.�q�`���˿�/�B�C8��+戽B\�����$�1_�U��mAV*�λn���h�����xg�օP�e�+��2yO6�&�m�k���mef��  ��IDAT�����ٽ��2L�X.�����}����Ii���	Y�]�Az��	����=�w��?�?��j�������5��_���_����?��G��?o�'������l[�G�«�/�k��n'����_���������?����?��������?�����/��/�/��O����ߴO|�����OlaA}��ƕ-�r�.��S�UF�#!�� @�\�[�7a�X���5���"�����>�/m�O�yJ�yÊM)��R�~�@�bۯ�������X��f�+��`�~Ap��6ķY��o&�`쭋�S,U|�>�b�W2���ӌ�F�	�!2� `��� =����WO��C~�`Mu�tIe)/x�����!�	��.��{���/Ʒd�R��֛�FO�2�z��ȋb�+�'	� `Q¤�c�P���i����G���;'.�d5��k�` L�6r���F3��%���p0NC����Z����h��*�����}~���Un��U��Qj�����Uf��kOӦ�J���XP+�'��7d*7-��T��%m��Q��Λ���{�=t�m���ޞ`]�u\bͺ:K�תX�%���-�a)/Ik]��i�c�B�4��ػ�n���m�S�d}�q�1�ؽ_c�9-���do<���$�'��6e��!��W�
t�����M?�E����r����>g'�fSL@��-��B�R���G�a�"a�,���sϿd��-�{1��b�Oi+J�"�̂҆0òP�T&���C!ÝI�<y�Q_f��|MK��}���b�g����Y���K �+�%M�=P����X7"<��
		�wD�]����o��4bV�'�������SmUl�A�&��?4!�M[�R�%3�����m�Đd��%�`v���K(�����X����a���cS�T���A�Pb���������S��;n����`�0��b� �*�-�<ܛ�(��V��j�U12d���/�e3�Y��>h�؏ڇ~�C����{�;�no}�[��o�>���������~����wٝw�n��퍎��-[l���6>1�L���b�ΜU�mYzA`-Lfl�Ot3�Bl�:5�lU������u҃.�8 �ڊ�|Y֙�BU8[V�f�;sņ-V:��H\��g��4�H`6�I	2	>ŕ�dE�f+�DV���$$�T�ތ���"EC�y�#��(!��*^�*Z�pl��K03��XE*�>��p�S�g9��DS�=3�h�vi�l3R��U[f�#)x
{�/��PAP4��-F�v9J9�g�,��V�ߊ��͕�.-��������+E�]h'�dJ1�B�)��8'�Jd�0���@ɽAD���B��҂`0�b������G:6=v���`Vw��+�<0����� �[��T��+.�M�����ޘ�,!��va�����(_:���8��K�3z�5��ﵡ���S�6Nضy;���m0����(�ٓ�z�Ǧ��[�\��;���}�Y5e|�s���*�@Ɇ���w�6۩|����A�љJr�[H��f��2�O���GmPm���]R�W��Cu� `����!JX�	o�W�T��#̴�~�ˀ8�ſ������`<����q�YXPֽ6<&KWn2ׯ�f�h���rQ
�	o�ko�*��1އ;�J̹�W*<���h��	&
�Y9qIA�P:�1��YC��q�&۶u�4_�~W�`����ũY++.���w���=�q�-���.*4�w���a��3���Jm�Qۣ�t�<���~����ZO<�:%li����X�x߽w۽w��4�N�A�l��]��3T`�P�[x��a���4�386H�e�R?aMPEΥ��c�N��|j�	����g�	<
�0�B(�ѡ�A{��o���;�m��������_ؿ��i�����/��?�_������{�՗dy���h^����y{C��췟�/~�6sqƶm�lw����v�~�G?���������ߴ�z���Ƽ}ᴈ���ي��h^x���eO�Ȃ^(�l��H$��C�2I`	�{d���V�$bj��Ĥ�G��G�D�b��+-��u�p����L��1.<�z�V.7U~K�CFY�[ˠ�'���;�2�RźbB�'k��㓲Q�2�y}�����h*�vzs��;��$�x����Z	[��Ѩ���ffmZ���vZ���)�s�$e�׫������c�7�-�6¥�Y��^��҈�B�c��K����^�E)]h MZՀ�b��[݄�b0��F��rfZ�ǫo�򌍀̼�o�6��&�\RH,�+,W�������j` ��r��V�?�z^u���,��#���7\\�߾hZW�=��#���K�����#�Y_�i�ٴ �KR�	%�?����Ci]�q��Z�;k�O��g��R�91�lq�n'�_3JG������;�X[����+6 �qrrXpe�rR��/"�<�G�@�(��]������&��3L���t���4n����(t�����?'eƻFu���-?���Lz}���|��]��|ɀ�6�`K/*�\^Zv�rXL��.<���c["N�V&�E�(�ּ���=L�PPmfaBD��.�(;�����=��y^0^�j�`���>$��Պbrss֖v<;�d�N����fٵ��Fp��k��{:�G�[��X��ڢ1�G��'후����ݝ�Q����OVZqY��ԅKn�$�=����FG�6?Weח���Ө`��#�E�q�W�CZ����]�+o\ju��MMϸPg��w�]������ʄ��uՆ�}rx�gi��0��:r�u;r�5�8}AL~�%�ff.ڙ�'���|����}R��]ۥ�b�蹬�5lذe�F{��v����Yw�	��D�+��K)c�;pX�&�a������$Tbz�\ȫ3�5v�P��6�n�ʺ+�R%���;(�2���^�k��U� UY�ǹ�}i�\R�6V�,]��i�ڒ�.z`k��,0u��At~]Q�f��^�I���paRw�P����;-��:�����J��uo��C����%*���Ċp����9��>w��>�f%�{�v<�K89�<D��{(����+�*e7�D�}�R�Y��b)�r&��|�.t%A�QE�"\0Bv� SLi�3ň! �HG�6l��2��z�	)m㘜���Z**�5��s�V��Ӕv�4㔬����Ɇ���by5Vk�����{��5�/��}g�~�����a�[�}p���GZ�gF�+��=�]�U��s�v�+_4��hYY`i�zJ�L�e%\��޷�[�-Lo������m�,NٳO}E�巅�0�~	�	��ן��%Y�̊R����`��]��b��պm۹�v��k+��D�Fsna���{侻��};-!k4��Y��`�K��H�z�1շ3;e/���wa�6�̒����5,|����������!x����LW�A��;u�G@~� 4�~ _�*"��"��,��Ꮄ���Ko��9}�m޶��G��8E�))=	1æ���l����R^U^�`��Nw�j����쀑LA�������%�gK0	��u���826 ���l�5??'M�aw�y�~�/�+U���E�KV�0�R��_z���/۲T��p������LT#��.�����f�0�q�3URQm��
lN�E�(=)�['���N7��{��4t�T�ZAL����§�����1���YS��#�g�l!�`Ƥfa��e1q �a��`V<�7c�����q�ȃu�X���N����_��.�K��v>�'xa%�lq勫��&�( ]�Q�̙SJ�l�Z����}᳟��z�����\�����}�gif�׶l��nbb��򃶬����*gHB�~fsv�t˦M���A9�h��m�0�A��Ev��-$�8�V�,�J� �UB�<s�V���{�������'a�'x��V^�d���,�ְ�aѸpn8�p:3?%x�����T$��WRfWK֩,���5Yy�e+(���9),F��baA�Y��.KY������d�J9Ooa��
�&>�֨X�^�3�f��j՗K�����L}Yx�*��t�#36�q�,UY�����~`w��s��p�f۱m��J�(Ĭ�ױ�:2����?#�u�d=�_/ p�+Q��ؼe�e�g�M�Y+�K�U����v��޵� q,R�Q� �KI�m�{n���$2 ��Tud�^����ꠔ�F"���+�5-�ۗ�ţvt�u���4�ʺ×����h�S&É��7m8�+%�js���wfiCt���O��+5L��&�k�&�Ϟq���K��#$��L�?�<p�ݸ�咲r%F�aU�1���ղ�PʆF�mxl�^=z�^z���ԹM`"d�a:x�R"�yG5���!�I�P�˪[��"��Pʚ��e[����nܭ�c�Ӫ� X
�\0	�M�l׭UX��6(bV?q�s�)���MB[�;���� 6���������n�B��D�R>:�u�
G�pu���V�Lq�Ų։YIL��L��Jh
�P��(�{�����C�t�vס,F�NKBd�{wCB�b�h�h� �%ƍ������~�l��-6=s��u�P�f��sⵄ]'L<@�%\�U��ۅ���5��^G��G�U)�ʯP�⨲9�́-�y�g������=r���	�*|QT���&���a	3]�L,b�K?�	*���"�����͗��F���>�R+����'�����!�Q8p�/�a�+�xy�%@RL��rp������mߞ=ʷ�^y�e[ZZ��;v��]�l�֭�k�vۺy��م��l��y[� �T�޶��%�0Q�0��24�=�ֲI�2M>�0�a���(�8��D5�����<�	]m���y)]���/)MKf���^O�j�Ĉ{�6J2eWH���p�8;��UT�p^��I�?��5��Xvm�ce��դ�k�K�\���%�����e����[����]����qk���]�`W�HxN�oK�)�ve�V�3R����u+�4sFBq^�@يKs�"��'Ōa�Q��oo��_XB�i�v���Z5���qU�0
>�ܥ��
Qބ�>1�q�;�	J��H޶L������m�q�e�VA���!��L�+I�]`<N�b�=�RO@��W�B�7/`	3�M�c�rz�ɝN���Z�� 3��M�.Z4����J����ׄ�#zW@��E����ҷe�0Q�d��pӆ��Һf���/I�H����]"�c��!��΃�vl�lk�¼�B��,�}� �L�~Y�)��+B�/~UZ��c�#��-!ZC}��Kʑq�}�.�X����?�~w���+J[C���
3���ͷ��n��]n�Z`��XYC�Q��F�\�K�I{.�l\�ʂ_6��~����Wn��Ƿ^�6�$����M�2̍�֘,i�R�z������엊�$^\(ؙ�R6V`D�X޴BA�pD<�"B%�D�R��5���H�0��7�%S������#����ݏ�`>}�yIB�$��D,Q���g=��
��J ���}/W��Xa#�e
{>?dI1��򟝽d�j�����?�N۹}D��`"� M8���pXP���>p�!��p�����d7��o�Ȕ�4�Z���K�3a_�� �u��7�/��øj9���W��KOBw��-�7ۍ7�`���B�pց��*nܕS�0@&������L��CEo �B����1f��h,I_A�C��Ҕܤ0�ö�r�86d�ނ6;�4m�}@�O�ި)mGVG�e]���H1��ɋo���;���O�?���?���f���~����!��Tl8�l�w�ه=d?��o�����z�a��a��V��|�6�v�����o����^�eϸ�H�hf���e	���w�o������?�;����߶������f�e:�q��~�?h�o���͟�9��?��;���,�^KI��-K7�+�.9�O�D>c#)Y���87cs3����81g�E!�a�A�% Q!�w\r��^Qr��슫���hK�a�cL֬�8뒷J�ؿk�x��+|秦��ρ�P�b��+��Ɇ2-�{��#�Ĺe�� Dg\B�#<�!.�^i�Y�-�nG���%Mq�.͠���p��������PZ.!�,C\f=bXL�f��n\������KS:�+�0TV����<��2Z��T]Y��P]�i��]�3��1x�0���)�p�e���V��j����j�2e܈�eh���y���}2o�=���Ŝ7[\e���8a�"2&W|�kOؓϽd��%��֑�
^�xF��bЬUj��ٲ�n��=v�-w��ԀQ���j	���kh»������ӱ�����)QbP<��\R��b�eeLn���Wտ=�����M1 A�˵[E��
�Yǎ ��L��5��,��,x��0t�2 "�N���wۦ~�j����z1��%XWfY�߸qLD� }�"����4�� 7Ll�V͢t���3�paW�؄2�����l�3�Szvy�#�4Nd�����Moi�J�d}R�o�aǏ���OXS�%�bغ�L�����?����\q�P��w����e_�.: ����0�QǺoIVu��7�lC��Է�r�ؗ"��eM�vx�}�G>hw޶ߖ�|<ș< v�T_�n��r�-��C�*/rCA��:�]D�����>c	x,������K����]�Y�*���^��Lس���߮o���K��/��^|U妭ި١�H��I�H��-�l|L�l��F�`X��;�:;�^����*�KeX�mT��w%)*l�Ђ��i1�o|�R������hhsKy�I~�}�/�zP����s�,�)�o}�zT_b�������y�}�F��>c˳�U߄��]��X��T�|�����f7߰�n�q�� X�q�.���u����&{��C�؃�أ�l�{���V{���������v����n�}�^{�#wIP�k�=r�����[��y�.{�m����iw޺��E�����l��;n?l����c7��i���v�M7ض-�.8�G+d������/C������,��--�[E�0�rR��$�]|�7���ȍ�.~�(F�yǮ,���Ϟ�y�%610�9�A���oߺA9���\�^<:ese�hrX���{v�XV=B'7�����BPe��"S0�&G�T���Ғ���Ôͨ����,���g�B�D�@$��9��/ش��-���u��F�U�u0|G��C��q�����w��!��Ǧ����U�6{��,��奝��k�SIHx��L��9��ҋ��߹m�M�؈�[Z*��:'F����O?c�b4IbU
AYnRZc2� �4"EfA!T��N�����e��]{������>nc#�62����a;w���K�C���L��ژ�U*d?N	k��vꕗ-!!; e����4bNQ�s�wy���`1D�º��|�<A�wFʂdf��Ԑ^)D����o�`㛶H�A0(�*W)��^��y�,�N�q$�,��C24u��[y��勘���{p����!D�q,2�j&Q@0O�s� ��O�ď��?�~1ZY�Ū--mf~�.�.��ܢ������W�X1E�����]����ǬlݶM���R�n�.���B�!cU��;������osP��#�Uo*�ƭ1�h���EDQ�����?��EgPh�����W����˯JA8)&��6.~��(�.�,�70� �|��ܽ{Ww�))ٲ���V��ٳv���S����-]����!�J	�2����}�*>ũa9�|�K�lU)N�h�'<��"_,(=�����i/x�EMH��?� ~��JR�ͧj��P��
�j^�}&��ނ�o����I��;��
G9�"#�Ǥ�wNF���wn�G��k����kVZ���e����:nl��A�ө��X�� z�B?��l˖aۺ�E�%���={�M�9!�x��8t`���6n������lZ�mT��Kxk��?�������i��3))&iY��P�#�1�-7ڨ���dE��u���(R�pτZ�f�#�?|�c�2bF߱��,���jG��O�o�KsS�*z���dH��>�W�b�W�u�Ru͞{��;�`��^ѹ�Y!;X�#��-#L��:niV��>����/��>��{������Cv��Ƚ;7ءv�}�{�= d.�>���RR�c�o9|����ϱ$�
�}�ʁ�8�&���T;];�"�+����� ���D���*��9�[j��(���~�g��1�0x���N8� Y9��Vw�s�U]9ޜC��[��Ԓ��ޜ����wX�[k���"������D��3^�e��Z��	�L���ȍ�ā�1� �<�+��7M8�y�� ���$����cD/Z�Qk\��(���º<r�/�����w�^�f�$��N*<p��[LX�e�e�T��	*�8Ѧ����@ٻ�$.eA'��X�a劕�@7���DkY5ԖlH�,�vگe���6m��+�Y

��?��v��C���Np�:#R�:�+� ��Յ嚶���D�~VF�Dc9|�«��8}"š�2��.��M���)[�R/��%2#�7Mʃ�ϰ߼%j��U�����e��E�F�l[
��kV�rA��&a,r��CBM���{�=�rɥ�����Vd��q�J�^
ς6(��j ���1�dÉe�U������FO_��zf�����)������	<��D�匹5�,qACe#�V�^���s�.�:y���B��Ya_�|aJ^M��ա��g�a��P�uҞ�}o޵o{��q�&�R*���d
<�y���wlZ�i�&-!���Eu5��(�:�]�j3jrȀ�iRQ@��gf���&yd�<%�j~�5%����Pv�Zg�]��gab|G����y�|�$gg�,yE&�L�m/I��l�O�3է��H�*pI@��4�Ѹ�<T�*��PrK/�*>F�|���Ƣ��NDba��
���TO<w�~ҝ'I��$k����geMʮ�}m|o]��|��"�U�eÛ^3��#)~%=�z��_͍#�|rSaP]"E��А(�yM�� |�(�T
��"�]��t^ӞdQ�ID�}���<��������&�Q	v!O�N6/0Ulc��'��c���켦ѓ��9���C�ϲ����,�G�v�8���,8��K��&��Ca��ЋC'�&��?�}�8u��石��P�q��NAe��E9D���H�'{0>:o�DJѯ~ă>�s�zĽ���?����C��697�3#��{-�j�֌�J8ڤp
y�h=Lb��ytQ�}�gހ���fl[ݍ^Z#�x�VI�7�V�T^GFo����� 46Ba"��_29q7iý��|$P"��!Y���3?�
�,�apBM
�[����lpvl�G��ۅ���A�hȃp[��{��vR�����H�%o����Q��Z�sTbu���QYM,.b|n���$�A�A�:3Jta��UX�~5��Q�X(�Q�s4�\sF��(�K[�F���S'-�[�Z�(�J)�2yWg/z��h=��+R����CB�U&w��I5�b�F��F�u��<r���	(!����M���*z��tAb��v���'@&L��T8K�y�.?��#�K�h|���odr#{τ���F��u��Q��Rx��0��%����ޓ�OS��$��~�7NMW-��(�>نe��\>G�k�֭�����E��r�&�9H�sb8)Aђ��
J�'E'k��S�4��ܛ|�� ��,x��$�_����}h¼�m�c���֮�.] �������{��nZ��{��^�X2� _V���,������H߫�Tp��V�P㿶��7�*AL��̑��]q�.5>��&`�������a���J�,�"�57��_��.��w踐�*F�}�){��e��ⳍ�jn!h)7m�}Χ�X	<�����G���:��"$� �T�H�ƾ��1�ر�����NA�ǳ� x�@�֮�"-����Veq���~T�e�+�Ut����J`-h��ŕS�=K;��@ez�._Çp��!��e�cgT�5�~��wZ�m�t�
��g���j�݅�R�<��f����!RJ<_0���#�dQ$���I�X��=���Tr�G�����ᱧ���Q�:��t͏Scs8|qϝ8���Ï<����cp������x��x���8x�<���ώ���>���NӲ>�#��[$�����".�L����x����i�u#�ưH�BS�Ә����U+�������f��g5�*/�@��ZyC|�N�[̂K@M�H���c�[����hD
�Vf�9��2y �׺@�%]JP���Q�>yGNَA��v>���b��ͤ�ʔ�G�M��l���(�7޺li����{e �����\��?�cs���&I�|1��T��)`6����x��;-K�sR2�_�,�D�g��@ipҚg��
S�9*4!A���)؄n��cx��'╻A-�:��N#I���՛~k�AJF
/Ϻ��k��i���P�g��g�&|zi�݇�kع��K��$2Ѳ"���D,!�0JA6�r-���"���Z��� �P`L�mU�>�nv^�^6x�֙Ln�5�(��L ֜Zr�X"4����)HX�,	I6[(��z�Q���-p:M�Ya�hi�M��K��1���Eb�Th�S������_U�5+�Fh��\�H�P�T�h- ��iqbs�����#(��I�Q*������z�~S�Z�9Y�z�^�2���a�,1
����ɳ�g�($l��eQ�S�������:�&,RLHOQ�cW�`ӦX�j�ږ�w�2�A�$�D�]�r����ݘ��r��yN�Z���8��Q��q>=Ъb4E�2w�R�mڰڬp��07;m.4)
�N�:����l*�6�]��B��L��k����ry+[�,wM� ��<����Sa{�xʃ觲^=4�������|�q����ގKRB��m<�?c�)�D�[Z��R
J �ںO��j ]g�}�ݩ�_|�M���	N������#g(�"� �X>+��O�^2���-C�IlD�zet_��w��TMU(�3|����LMN�B:R&�@0�G�h�(	_K��cK[�Ux��E�Iŷ�J��Ȩ����֭��uz��Cattu���o�6�(𩸏\��/!$!G�5���K���iJ��4X<NkKQ��(�_��5��vm[��.���}]�׾�c|���ȉ�8z�2|b?}�<I���3Tr������;;�S4N�H�v���!*�c'/���c'.����a=�;��'�D_�����N�38|�4��p{�����3��i�^��#�x�<��a<�̳F��v^��ľ�� R����Rx�)����/��5-p�yݼ��Az�����O�)���Jف򌆳D76A�'��@1іv���@�����V��xx㦭��肋����+�8C ���Q��}�:�E�*EQ�,�Ls[�e"%�j��M�	��z>�W��߳�"���*�i��w���w����9~����ۯ��>����݇�~�q� 2��o!l�h5�$�Tc���rGX��]����.o*ok��^���o�F$-*�C����+���݈={�a��^�]ǎ��X?B�WD��O�hkX9����=��#B������Q��\v�Ѽ.��)�7�C��߉\9Kᔳ`Om�:}QZ�dB/Qi`	�J�RW���>����f2yZ�,7U�'���A�2eZw�X��� \D�m~/<D�.}R)rV��˴4��V�Da-�j��ݎ�b�EʩFE*Q)��{�Z���c����⩯��\���?�c<��o��c?A��QxKE�%��ɽӐ@Ц�ii{�>i�(��B6팹4	
��6-���Yu��8_@g�

���/��/$���=�@AD��#����Uz��)r�(W`+��?�g	,Z�D�B���V`�K���4�,&l	uё~k�A�JA<O�HXY94�}�u��'�����?A�/h�B��4ꔀ�|�<EH����])���)�+�z�[�I�X%��$�8�yM�הk�2��X>�e�L@�:�q�j�~��×>�Ox���d��B���V�,[���"	���V�2kx	@��Lq�6XG��ж���eQ;I~��r6�^�Z~��7�qvGΝ�s����N��w���@��g)�@���,����J�{��w��{���~�7�@%/kM���,��&09!p������\7ZV�\�rc��j���X�]�֧=�]&|�F��>�Q��QkO�y^��r\���ۣ^���2a��F13O%-�4����s��U�y�z^ �A4��hb!W��O�#�n��T��}�m�AzWf��މxr���,I�A��p?��k�ٳ���\	�j7jM�v&Hv��<;��r��G�}p�b,g�P��
!Cp2=�ƙs�0MKZ��j�v�\��đ��b�,�K���@d;���&u	���J5���6ߑOic{7H�m�VTb
���O�y`���Z�k3���:-�O2�����Rڵ����u��n�
����+� %��iR��}$D?����EF�=�v,N��<Q�}��!>����??�o�>\�2K�#z����Q�����ƷB�q�(�A�ri0R�<�XA)>1�1�>�3?�Qg���eYz���.,�����&�S�Ee/��6�0�P؅�I��e��$P*��?��T�J�q�U��n��qM������;v"��E���@0U�c^�m�m�b��u�|�Ļ;��yq��M*E��z[��BI*w��`�,�hW�D�S�y�;r�Ǒ�gq��)(P"�`��h�D܆�tQ-#@�I��Y�|�<��2��E$�&p��+�V[�6)-#�?n�����i�{�)\x~�����E�VB��-,�4v�/<��c������`h7��rtq�NszE�,_�[���w�ƌ5.��F����$�4os��&�I�ʞ��L`{*}��&q��iLN-�8�w)e��{m�r��4�����O�߱V���^.Q��I�ٽ&�EK|�	=���3,G�ډ.f��S����"n�z�|��w�}�kX��ҋ�������]��2��x��9)Zk��]�x\{�B^Jgbl�2w�"!�tV��_����Y"-+*cMւ�
Ek�H��µ�-ׯUGmv�e����uj)0<���.^�u���՛�hw���i\��3h�Qh�I��{�Q
g�������I���e4²/,��"A�Z�
��H���H'������|
gϞ�U��ԢM8.Q�I�I�)
\K:I1j)))=���P�G.c��(&&&��3{i՝��B�x��������[��~)d,Ë>5}a��*�f���iE����T�*/-��d,��{A�.|n�2�%�0�e=�H������߻�C,G|�2�LO/b�
���'HYn������g�y)�ې�FS*���wj�t�357�A1�����"������A=TŘ&��X�f%�c��(�����<u��-hױ�qK���v��O����9�u��|�vm
R�p	�VNy�	zY��M�"��ʨ���5��<8�e)��X2����4�S,�Q���5��LRx�k�^w�;����=��������P��Mt!���By�D��5��Y
��������PYx�ܩ��HT�J`�6i���ov��]}J�E��,5�KG�wnbbcd)
)cnq���[��gH(���"[?�&�������k�&�Q�r�lز�(�ft�HϬ,:�(t6�æ���ڷ��vnE�#f�E��%B��*�bT�2�&h�I��-�v��z��FTTd�S�����Cx�g��|��ַ��#����}�A2�$;R�թr�z�hP�B��B��j\�"��q�7���@ͮL�rIY|�;�ۮ��V� �r�(��E��#�A/5���A�k	�l���Z�=g�Gz��H!
X7A���)/nz����,r�h���K(泈S���FG�B��F�uP����"�U"���u�Jc�,���38}n�\���H���� �����,H1���$��R���XD��RzW+'l��4��zh�,e���/r'֪%ZTZZ_��[������s?��������b{���a�Z��e���ҀhV��&�J��u^��&��h�_GZ�ş{���>�����Ď-�y܉Lu��K��$s���36ޢ�8��QRjyQt���2g�uN�2�>f�u-D��������9��������i9rZ0m�KE��F���	���Mz� ��BT��T=�4991nA�\zy>a�
���dD���c������%W*���ʣ�d�,�)?������6�mo{y������o��ߎD2���YS���i�^���ED���z^I�Z���HN>%_�4?�%�#B���rR�S1*�1AROW ���"ʐ~��̙�����ź�뱊�ך��uE�V	�kU�ek򾋆��}.���iMY�ߢf�FcQZ�1�Ϝ1}?etX�8Be�F ���T�%͠k֭�����e��(9k|�������֢燔޲r�<�5`Қ����n
O��L�����ԧt��j]|!��R�7G>��/�O
���F�<GP��ʎ��lѲ�c��;�*�y�=��\¥�<��>�X���1@ȗ�Y�`W[7��}$�2�{v/N��L¢����d\1�!�F^�OQ�P�PxhR�U4E�DA`�
&�����I(5��LX:5+&%���|[��m�L.d_b�OI@�z���c�'$���hҴNR`���1~�i�
��{uٹs��Hn�-{�å��p��I�*�n���?����[��߅l���D��*3%lڲ��~4o���Y��I�" Q&Am�8�	���$���l+
;�E�\.�
�(u-d�U����u2�ؕLMO� *dg�S�E��D��2�溺/V�\'A��@l�:dKz��mge�p�����"R����!v{z�
�>�$���m����f)OKh��"6	�F��]C�%�=�>�v��@�TFvs����eI)(��6"ѢS0HgN��s��y�:,�)bn�`���k�o�_1�
�2v�藺�pW��'�X��v"������E���Rn�YC�On|���[���bf�d-�*M�]�*�c|cng(�MH&���̽�eeI��n2��-�p�M;���k�k�lܰ�揉:���R[I��2i{�E�Q�)k��Mo7V�ZA%��{����/}�y�p;�9�Ӊ�������v��D@LeN��u��Z�'!U���
��gA����:V H�����ďj/]�OM��-��́�ƫI+�r+��U<��^�䁧Piz�a�6ܴ\�	c}|ZB��_;ԋ�w��X��
�f2ʙ��.�f�K��~�f�)�wRQuDH��	}6}�L>��� �lѦ`#ɣ0�q=���o��xO�m�n�w�-T�[l\���K�3Tq�#=�d��rT����)<��	�!�>��ܜTzC]�x�L�)K �����<�;:�f�0&Gϣ��Pw��0�Ͷ sH.��p� 0Ypd�wp���)���c��3�8B 0G�VFWw����+=�PЍ0�Q�Σ^�s/�T�Z��T��4��K_I���y�$~K>�%�j�r�{y�4������׭���x��[S�d�HVʺ�����8�^�X����h�e(l�?@,�B1��ۭj|%�L@O
�\ݒ#��X,f:F4)�.��a���-��a�p�2u<w|c���� �wnض+(gH��{F5�vՖ/��)����g���������_�?��_��|䗉n�X��2��ȳ3�\>�gH���,�J��Ae��TcY��ML��AR��F������q��*�P��8�K��-�!0^/A͆K���E`.��gR6��q�'� �+�Ʉ�<�Ʉ,?��RYD�I&t��Fu��֮S�����E��2D�
sO�i������[��hQiٔ�HK.i��J��%-��(��u,��Á
�O`�8��+H�{	j�dp���Ճ�f%�4���P+����Z�ٖ����mw�Y�Ѷ87O�@�Ë4UĮ%!kBq�vц��'�QTS�C5�C�G�W[��TY�ʣM�ah���2�%*��,ۗ�uiI����l/�j�(��+F�\��o��Y&�'O����k&܌X$%8(�i�'�����	 @�Rr����D�Rb8NM�H:j��Ġ��mc�|���+���jM��Z�iS�kV������W����������>����G�?����������������o|�O}���'�������k�~�Mرu��~�v���v��X>![�SEUk��������@C�]ª�z��-�����뜔�\�R&R�/�S~_������]�Ȝ>s<�(-���$���a����H1,��}ܰu�rY�A�v�8�)W��i�MP��L1�슪����;L�9�$M)C9���,:��&a�y��pe��c'����uQ)IFttv�om��M`A
_AzuM ��$��&f��yZn�mT
�DK_i�V_��y�����CqZ2:$���R4�ŷM��LV���"�(��n���,J@W,g(�`s'W��ޤ��8��'I����/��iJ�ʥHQ:��w�2��"	�G��o�wщ���^�9��`D�J �yݵ��_�0�N+���y��Pj7͵�'���ϊ���Ib"}��W���!�Ck���<8��d��(c�����.Vd���S���D��A�y5c}�
-���:M�#G��bS�� V��A'�y(�3��y4�7�Ɗ����kq�ݷa�֍�����eC��#[���꡹�c�V�� ����Y!U��R"*����b�����q�Ơ`d�m@��R�91�����+5}�䈶b
3���6⚵]6��Lz2ѹs��&CQ����@sհi�:["cߡS8~v����c��m$R��K�)I��4h�>��w97Oa�����8L�
ɍ�ᕈG�<��5]�T�5Zl��V; hH൷]�AZ�񈗊�B��a��I(M[���j�;3�~�S��_���7���M���F� ��O��5�E��ˮ��r13�P�_9s�
l���R#Ӓ�%� ��%�8;��
����v!>@e��icj
a6+�/�K�n�\�2ض9A��Ǿ�!���v��Z}\L�����5�%E�C��Q�d�ɨe2��4Š�ݻw��W��H�(�S��r��V��)0E�ASZ,�W�6�k���u��:+��V��61�,�V�N5�%_&�3W)�
�y��"ѦM���ܚU�X���֮�+q�-7�֛����+{�b���	���ȃ%ZPZNcW��ƃ����:�D-��R�^*��T�o���R�RZ�CkW��[��x|���H�;c�����Y{���R����.P��mirj����G�@ָ>|�\*
;O�D��%�aUO��Y���[�q	�<��^�S9S7�|-�y�)k<���H$���i&� P$!��\���U������jBt��"<�R�l���D��y<��Cp�v�zlٺ]]�6���u�>w?y�� ��*o/<~y�ʴv�:.T��B^�4yܴ$X:5�lj� ^{�ʹ�YVZ)G'��S��̅IT�8%�Ba5`�z��ҝm�M�H�ٳ���ߥ�RT�Z\	�5'Oc{Č�ݖ�#M�IX^5�r��~��;lL����R:��v�ډɱ)x��Ǖ/�ѮM��r;�6]��Z���9{v������	w`��MNR���^;w\Gx7�y�f�\��l�L�-�CʌO�3��B�|���cX�"Z6l����ȕڰ��%��Sֲ�Z��_��>N
��P �	daH�H3K �V٠��QRH��s_�c����&d���ç��w�'���#~�֯��=x߻�Ň���Gރ�n��B���Gs���۲7�.�c�A=�o�Ժ��|�~�^�K��)bj~���1E���h�W�G_� :��l���ʱlm֭�ee� �LE�}��uS��cT0^$"!�"At&���$(�4`M�Q���(�&J��������/�Cjv��@;6�[�7��F��og[������Ƶ�d�W'�wߎ=׮�*�+���7��+��v�B�f"����K.
���"s�G�̋J��qvml)A�קB�5���j3���4�_5b�ʼ�am)L�y�?�wGr�S�K�k@���w{��[�R�D��+�єl{:�%����|���n�h
Q�)]\�U�b�ƅ�
6��ɽ{��A+h':����WolSf�T)SsWr7$�6R������Ru��\)B��@�������J�ȵ*Ԯy���T�.D#��\%�׼��i���	���\���������i���Ts%�4KZbt	�H���GE�w/��Y�r|!B���c��e��*�v)��wyutܶe�p�L�º�~	-�6h!}	#���M�P,���SO��g��P���q;Ai�G�r�rR��g�M��|ߺ��'�"�ʸ�������1=e��#ظi��B�Lv��
�q@��Q��]z�zi�u����2Ҵ�˚[���b�J�H;��)�Z��e&���!����!EXQ�	˨�U�UX�15�Fe��P.мD��UH_u^�o,a��S��b]�����Q�	nK7��&FgӶ�j����-}SZ��$@�<��԰ q���"�Ũ��Ж�>5>������.���Td^�]Ez{l�VYS��(��a���5�C
Q�v�;�v��ٮ�T��ӛ�� �U� ���������?�\b҂�4����{z���AI6�������p�-�{��7�0�F�g7֮Y��6��`�+zӦ״<2�F}&��W���5K�Ⱥ�"M��E�Txl*<�.,e'M-t$e��r�Q5�gK<����\?~�q|󻏋P)*�8�o1=>B�6ᷰPFz���N֭^A�W0�o���D�2z����b���?m����cyH�V/�uIh5����-J��#�)T��=�]���D��|Gw?��d�	>ărQn-�4Q���-�2
B�lh	 	��V&5��X�=r5��=:� ���uL�Ob��W���׆P0�D4AF��(�578�`y�|f������H��v|��i�
t��O��Q8s������S�]ݦR ���m$p�~��	t��(L�L�	X��ɝ�tmZ�Mn��1[��H8(	�Ġ��*�����uN)��T�
��S�	��X�c�D�*��E����&8�4�?`{�-Y�������G1zy��nC6/Fe��"��8;�����T4멜��K�zb�㚶�M��|���XJ�,�" ���ԥ�+*O@Om#�_Y+4��F4"TXZ�D�o��S��ss������Z}Ds�4�@���䔹^m"Z�34n�^���*��)21��Y�Kt�k^���V�p��.%a�'K���*|��$��B�-\/�'f������4��"��P�r%�!�)��S4��i\~��\s+���MB���Ȥs���KT��?��V4��E�Ϝ9K�`��+��8y�$��Ƭ�.]���G��i*߇z���~|��_�?��?�{��.�=����)*�%�W#����K����'����](%�-�Ru�(��B[R��B�s'���PcI'�,����J�
�����)���A��%,K�/����yJ��8��Ҕ�EZ/W�@�~w��FcI�	wK�X�S�/�+�o�|By%f��w5�`;e��
�˝�.�R���}$��5��d�g�
r*��P�[tyY�	j7���1Z��W�r�f�-�\�U�q)���~���(fӤ��Y�rO���L�-o-nm�u��5W`ݔ?�J~��w������r�#2�{�".N��@�ȴP�YP�� Ӌ�\[?��+q��q~~/N;���~�˗������<��;z
G�����><��4�+���Dtv���4_�Lt���۷ �X����J�oX�*��A�6���eE�B^
�vLg��"�*hE*�,G���Qz��R��cmW�c��n,}f(�3u�
u
�2(��At�T�J�������8�T��SYN.�;��˗�ä�5*�u Ǯ����EKP�Q!��Ԛ+���2i--��o`blǏ�����Q��j��h�ţmx�{�M��³�����$�������#�S��v��6G��=8=UD����X�	�
j��ӎ�����vu����c4���\�U��Dea��DR���wC��ٞ��w�@cV��h-�x��7"��E��,�-nz?D�R:Q�d�Ϟ:���.�TlC2ց����A�\�EZ�O�-�R�|a��}C}���(e琛��������`˖�D�Ic�;)
VL���xؠ����\BZAo��5 &F�����ϋ�K�I��++PL���X'K�F�N�'���]��xR�Yb~����w)GES�z�ޥ� ���lT0�	O*3��p�b~	K;����dep��;)��Eiմ�\�"S�h�O	&��ή6�B�1JY�Ԯ�W���1"a�?��CI�A�^$�m�<�b����o��?u��Yɡ	~���"� � �P��?��F�
,�p�����#�y�������F��S)�l��/HK���y_�◨����c'p��i<þ׸܅��_ym�>�#ǎ�
�s���C/����W��OPA��-7_�M�AZ&���8z�(�^�h��w�u�z;m�7���ϟǁ��_�qѲ����0A�"��Y�ظ�w�`��κ�<5��Q\�}n�n����~衧�ΕLt��51�)Q�7�7qh0��(?�l3%p�����,���Ӻ�M*(E�*�P��B.c7�.���gH��mWg�������\��TJ�JƢ����9�N�:J�!�� ���?��4�I�ru�DKԣ�c)"������0AiW7���-t-�F대Ц�P��x�mw��9֙	iPQ�eM����\L��Q�j�?�\��Ztwua��l���k�4���wmB�^����t2i���������\��؈��y[�p��n��tu��ۣ �Ux�ވ��}l� �����ܓ{��}���x���Yx��z}.D�A
��ci��d���ŬRvb&);1������Z@�� �7�;�b���������W�O��-|�?�C��SϞ��\�
�M%�G:_�\����F���W������5H�V��p��q<���x���05:��5���3$�4-���y>c�ż���_�l�k07��g�~G^8d�w)ٳ��yVN����3s3Dլ��<Nb�<#)�*k��x����dH�$� �E-��$�9
��7���P�1[4�a�4$;;���A��9_�nPq� .3����Y�b�Z�`,��t�V���I̒�(*����a��$���K�R6����x�H�dj�V�(kctr���	 �Ŀ�y5��8bn�@�� �&�
(��-�7�ZV�29(�H�#kM������ax�NW�J��R���"QD�6-�IVE�:�U�,�`��O0�D��f-���B\�Ԑ�!g��	I�_+���O�F�5�{�I�G�K�NS.A�hH9�ʫwh�������vYs���2�Ts�Y-7���@�~
M/k0�~�����R��]�X��D��MI��oؓ�|hɐם�$j�ZH�"vY"�j��.:イ��� ���ʛ�[@����L6���qK���Q������(������o���1H�6�$]kr���4<���G�L�Å��Ē��m� d!��rYB�@�y"��`h�Z$�V��j�Bn�� ���7L�כ��,[�7?;#��h�X��j���[ļVT�����ڕ�YJ��O�%�(g�Y���a'lXD���M�p/Q�P�*hIѧ4zxLK�Γ�N�I M�
�'�"���'H{��&�m�8�P?�4�Lq�_D��AM���m��5��n�{ѿ�B.iџ�^�"��W)\?���)w���"�(������L�%�i���!Hn�	*φ����q��+�D��+�J���HmB�b$=�O�zɬlkv�A>����}������o�����>�ǿ�{������Kx�[߈7������?���O��O|���g��#|�?�{^wQu�Ec��c%`$h,BSۋ%[��|����bۘ`u>%��AdK���B��R���8G�YPFZp�4���Ri1j��0:��ah�l�r��*���q�Ә��R�i�x����&�H�i��8~�y[��D9d3e2��3D�v�}�#�N��S��Q���8�g?؄I��'��u��4ت�M
%��r-�ش������V�Q	e�$� ��\�o�[��L�/�FK/�z�ӺH��M�hkg�5)Ī�ddZ�f����rA���׭C�h�B���l�Y$
�Rh܅���;����CTe* ���{���H����4ٝ�٠U�ݿ�^�Uv�;g�-�ÇN��ߺ��P�R/YĦ��*�e��f����)^
bÈ'd���^����t�@����i����������4�.�'��8���2E���o=K呕�]
���P��y�n~jk�W�:�$��_k�"o]c�rUt̎/��]n;�/�p�6jݴ��]R��r��*�B�Lk�2��Sye��qT�|�{(��ko��D=)��kS���|���#xQ�ub'��J��Ւ?�
(���t%��$/���b�w����_�;��[��?�3���?������?�i���o��ݻM�i2��Hm�I���s�_��K�d���Uhc�k%-��ܒ7�6�� �� �1�a��w%��V��� �YB�׆ގ0U=�yv��k�L!zQAG؇M+�V���r�R)\�ܨ�<KT��`���^͒7
����n����y���i'Pq�w��]J�?(_d�����]r��Z�j�Q���(�%�]�=�]˷4�7�&�&-
J�I����v��D�4%DQ�D��������I�	���5�K:�鹢y�p����[BZl�fp��uB��gh��%�V����y��j�����JA���|׋^�%!�kTtu�\^� B��ϼz�]ش6½���H|�d�,�m��Χ	���ݗĪ�}��7�W~�C��/�׈KkL	��\0*�����U����{�]=�s����K��~x��G���<�%�,�3JA؇Pt�W���=���y?��]�~�ݸ�{��׼o~��p�7a�M��"(�Ȧ������3�6�� E��hү��������:x
O<�,F΍Sy�}#�����/*�=I�*��H����� ����2#�pQq�y�-?@�@�F�� ���?e.QU4�I%��]x�o����l�6,(b4G��3D�Ju%¡e�F�
T6�5�1���*���u�Ԫ^�&
p�&X$�{{�v�Pi)�+r��b։#�A��9Q�|!?�6�^���>m'Ôp��$�|�kv��6���f�����>�Gz���fɝc12�VY#��b؜L-�i�|�)=y�(�pƘ~z�x�,T1��RHT�8Jyṁu�2�դ�r)H́R�g�O�Mi�=GǔE�V���Vx*�ʤ����A�/�vk�je�M��l}:�8�i�W+T��k�skW�G�p���C��F��2�O>�U�'	�
���o���3��lJMҤ/O8	W�
� N�M���4ƤOYN��^���<������=װ-A+M�S"����_jͩ����Y�2d���}��/�ʯ��}>���Ǜ�r�~�밆 L�ٶ�;�;a�h�i�dD��K��"�.tt��|n�/���Q0���k<!��M��c�M��D^'��:�~*�
�|�HP�k�T�5��N�ҡ�z�JF�y���}f�I1�h嶎ɫ֘/�Q�YEt&�T����7]5*@*`%����� Pc9j�<iHѝ�@�I�qbQH��W6ޒ��#�o�沶� M:�Jޭ{xR�&���켼P-����-p���+(֭ۀK�G	4�0��Ņ,J|�y1���Էr�;�!��~����Azı�t~Ɇ<�[��C�6�����z����h��)`��\>P��>e� B��׬�J�BuP��k1�D)��e4���+x���Y�,�ّI<��0~��~<��i�r���}DJ���ɈR�b��&.� *�Ї�?m��I�-����1�Mϳq.6��!B
(z�N�kHx�٠I��Y�z�+��r��ٵ+Wl�%7���7a��mعm�������V��Z����َA��>1>a�Sp��8,,022�sgF06:�Φp�R���GQb����N��B~*5*�z��^ō���K�r�/�e��� �'���i�QR�h���_�A�6	��xqg��]^��m"tч�Ր)��`ڴ	��>TIX9�_�(=M�Z	+�W�e��"��5k�����E�))�yk��ٖy�^���0��N����)c�B�dKݰو�)�x��倱��P�\�힠�];{a��D��Nl�~ۤ_�\�<�����y���9�`�\��6�+��elN���*���h��-a�j��Q|2�T+�E��%
e
����`=G�,BKY+���\nP)U	F1ˍh�P��f�I�)��!�}❖�#~p>�g�m�O�[����׻~j�"�бO��м�㕛�*OP@;���(���>��f�R��K�&�~�#�ɥ��~�3ҋ�;��l�o*=�}�=-�
A)�!��.%&�V@�8���Ш�	S���ʬ�)z���x�'�3��~�7��'�ۿ������>��O᳟�,~���ʘ6�S�I���Z$_�8uG�� Ha{�؛,�� @_<!�}���|��M�ȢLeXQ�~E��b�N�^�#ߡ�<KN�V�R[�����arz�/\2��dg�Q���E늚��@�ʇʰ��@,e�( j�0E�f.P%r�G��`��@8�`Jy�˝��ߢ�Y*�6
y�b)�(4&�
F�U��Z��
���=/�������/��A:��M`LNM���bR�hX�jVz0L��d9�Ȥ��Ej��DE�8͚_�eۖ啦���j�*k��T~�N���Wۺ����Wkoey�O�<�+�D�D~혟���i��������X���l���$����>�<��O�����?yO<} {�>�XR���`�'�؋'�|aZ���Uv����}���Ht�����R�Aܭz�O�/��oD"�d���)��4�A�#��I�<��l�����%�)<J�Ȏ�c����Y9��6�L�m� �V.QWOG}�t�;;le��gO}�i	��w��+	����<������GZ�Mc��8&�)t��@Z�0��*l�B6�8�o���Xye[�.�Xd�Ԁr��ə.��cb�H�܋�;�t��
Q�G�� ۍ�
c��T�x��x;���$ ���ƶ�]�g�4>�da�j�_�l<-7E�*Sz��ZkVi����g��${нf=6�|'��}H�}�xz��H�*�&�v�QcܛUַ�N�e<���m�ܢ��5r�h�a�B�IK���fA���D�Kf��n�n�p�Y��V��u�������re7�іd6�#�k�eI�)�	��B�lM�-�R�#	�`���7D�E���t�%=S��pZ��U��y-����]�uvn�Nt�w�?)-Y�΅�l�֔
�R�N���=��C�YJA�L p3�?�#���ft��i^�m4�\
M֥+m��ˬs��}�̾����g��,�����O�O��w�ߩ9h[H�}�+\e�X�u+�q��k�$J�Hg��<9��	�)�^�e�:�?w�ƅR�Eʋ*�V^i�ʕQ�\�ɓ�i),�Е<����c�é)̑�eE����]1���+p�2B˓���
㷼�Z{�Yw-����:?�@���B���
9,��Y^��t��$ Rf������!]+Q�׷�|=�t�x�Б�8p��f�ȗ��H��mM�(QfU�em�VS�p���Q.dH���!�� I$��B17G;��I�>y\Sc��f��jI��z��M4�EJR��W7�\�^�����ٱ(�ڹxD4$e�͢1��#�&��'� �3
bpx�J�
��5@;�Q@�V���Z�@��~����frf� h�Ɠ��T]lCy8�T�m��c�Y�b��ʕ���=h2i��Y �d�%c~�y�th]��ǩ�X��r<}�5K	��bnzAV�]Q@�E��\s�v�!�iu��N��#G�Ta�k�.�)�)�4P�b�0v��l�8
S~j�!�Bδ�䄬x�Uf�έHv�m~�\�r�Hص&���[(���12�)<"i�5ϰ��J$2Q�*�'��2�	��d
h�i:��P�F,*�ʎh,#!&͟�j>��Kgq��Kh�٩|/;Gcu�=�4�3�D�W���*O�V�/�Pb�<T�~_������A-��bvo݊54�{::0���C���qz(<�M��s�f+�b%�$�t�R�E�ϹBFSEt�߉�k��-I-��K�#u��SDrèn"$-IZ2����W�ƺ���M�EFt!�;�ލ��e�M�y��X�b̑9����M8'��-6����b8��\+f��/j
\�8B]���1$DD+����%W��x�B��jT��4	��D`����N
��%g��%�s3ƨC��ٖ�x�|*�Ή15֪�[�Xo;�M4��uƵ�)�%f�oS���eul����^�3M8�)
�R|z����ǔ�w��s��h~���|��j��Atj��նR��ߞ����[���O�t��j�������Otl;(]�#Ţ1EI���� ���y ��/"�g]T"K~�� jn��s{P��b;"m���X����hOw"�=׬DG���eZ�ן��I���G�۰�_DAj*�@�V3��(����x�ϼ?���� ��w��o��.�����[��V��%�V{Z��!�
�@��}�Fg�Y�I�w��5�LVy������Ȱ^qs���P��KT�%����ҧu�a��"ŅI�Җ-���f[Jjn��E8r�'	f�	QZ��U*^-$+ŧq萿�[�߀7��v��]o������k�N%�۝�A2��k�q��x��ނ�8e��I��EE1޲��0E_�~MMӧ�zJ��㗶�2A|7n��\�|gO�z��Dö��{���*���_�䩐�Co^���v����h'�ԂԨ�d}	�j���.���4U,Q�R��T6ʅh8jt#�[��E��+	n:12���N^���vJ�xwݰ~���«�3�u<��IL�눐Hl���������,�پ�ܺ���x���1=[@(��!ڥ�u�5��������m��X��{�(;�
BL�u2���֝[�쎘�&����Ov�����͎�A	�$����,�i��L-�G��&��<�B��D���N��0͟J��z�@�I�טD��N�
�eRZ�}rr�V$zʈ%�1�HL	Z�o�(�}����Ķ�PhA�x�֤�D��b�c��0n��F۸U�D>�e��$�0��	Z�[v^�]7܆��uTx���1?� SҒ*,��A�K�b�+39�h��v�lX���2�H��/o@gn���Xm)E����m����(Y�L�$�H"l�-�	l��&oی�M���D��#�Te͑8)���o�&�Rx
���3�P%�9x�G�W�c�ּ�
��B�x�1�akm)�W�v����y�� ׼�M���E����ϟ5a����Rz�2vg?�x#�.��Z�^�2V��y��,*|�"��x�R�dk|Ц P)0K֝����tLm��֧���ڈ�OnΧ�p�-lr���Z/�9�qF1��R*���js�_�z������c�Z����7R�ˇ�j+EJ��K�.*k|���g���O�H���C�^��֠u���wjF�L��~�bUk�Q���w�ȡJ������I`��#���k_�-���2�K.����0��6TĬ�Ҥ�|����|�	<��98p j*�K�\�;v`�޽���3�,`"ZR1wvw��h��tY������a�����z��_A�V�7څ2��3(ZU��A��3+u��'K�9�.�bDoሗ ��=4��X�sO���x�X&>W�m~*U͕#�f�e�+��>�������*�>l^?�m[��m�q������B܍�o���^�-лv_c�ؾ�-w��o���ה���ٷ�f8t�@$/��Ϧ���YC�{�-7`��%�=}�����iG�/+Z�xFֶ�Ј�R���L�kN�ؕ1�g�[ē�/^�U���T
S:v�"Ƨ�_�y��E�B�E�ʛ!��]� aQ�=شi+zVF��p��L.�R��tFp��k����66����K�+�L����H��������H��ٕ:�9�<����v��Wc8�K�IXF#4]i�1�ɤ!e)"1�K�Ӑ�_6�j��A������,�pr��~�q6�4��4ff�͌�&�EQ!/6�dr�h� �\,��i>�d\��}�m������7���'"H�S��i���a^�����ȥ���:�b`�~�^���p��i\8wc��kD�}X�a;�mٍ����R��6v��G0����E���s��t��)у��5dZ�!	��K[��[�^�T�~i��P��EPI�2����4x�g`�H92��BE�K�D�T�l{efQ�Ȩ�P���by=��Sɺ��4?M~~-����M҉ܺ�ԼM�V��ԥ��A R�ϠQZD�^�"��P-���b��ظc'��$J���@�Zo�}?y�>���\,�r3r��[��h��/�F����%d��חS{�zm����Ρy��G旒3��v���FZ�S���-XkrwY����W�%�&1��>u~���]{K�i3 H>Vyt���u���V��{�)a$�k�_�j�QsF�nRQ�5K�~჏�g��_aj.k��B:��#hx�i$�v�*iEK�	 ��2��i�cR�F�������B�=�����_������{��E:�TC*���_���Yqb�\]]]����
ZCCCƣڕ`Z��R�����i_�ƾQj��vB�$Μ��������{���$�r,;���� �Y��'&�h���T�<F���'K�aI�V|��ExJD����
��#��s���s����)O�����N@W1>:������-�3� ��baj�2�2�Ŝ�ȅ��
۶��!�g�C�75@�����Eu�nz{�؞�J	�:�E�͡��h0���z�40a��s]]�6^������U|Q�����_��+��/|������'Ϟ1o�"����5s�
8�K"`&���E�<&Z��ij�ջU�P��c߸�
�\�{�岌�I�B>+W'-�=���5��w�y3\�p���K�����֮�{�Pȷ�Ab�U�9=Br�i�EĢr�8^ڝ2����ݦ�yi�#����i�,���bͦ��,
^8{�.ax��ҟa�g(�R<���k�T_o:��๬&]J�����U%T'�G�v�jy�����L-7��\�p�6n�� f��)�D*aZuQ���c���X�q֬ߌ���DN�Thu�>?�����dy\$GE�M1Ҡ�j`p�&${:(�J�D�K���۫79���
���Q�EPc�����k�\�"�H���4��@��D�
RjPy�lSa�%�^���E���MK(�J+gP/�in��@눇�����0�jq�H0�>��bߌNM��+$���ۦF��E�k�w��#|��?���<��r���r��<�H�r�h.��F���7� �RO�&�#�kK������7	c�M�U�Y�Zl��	E5��))*	���٬SA�M�-r1�*�����?	YkSY���.���զFqF��d?	���4�%�I��N��b�M�W�S�(pC�̑���?���s��+�)*�H����&m�C�Vy����۲@�0O�8IY �f��`���
���s��������I�ņ�ۑ褀�;�>��-�"0�qR	n)+���M��y�x��ކ�w`׮]��Q���/�_��	d)xk#����fYI�V��
%��6�o>�=�ٿ�~�0��$<Tv�^�%OZ��cK��Zz�����m�{JD�14�6M˴Fk6HES�"��,�j�H���R�g�T@������^$�K�X������A�QZÐ��t"�H����+��zE/�:�𳽔�Z�ٗ/_tܚ"�^(����I�f�}��G���EW"�Wn<x��|o
�����D�\�2��9� ���䤭����iLLO��%Zw&�5g/��*�����N��mܜ,h@��ԯBS�Zi�ч��^�kͰ�]���r����3<��)�dh"�:�(h��R 	�uP����;N+σ��nK���D(DU$n*V>��p����w�q-~.RH?Fd}��-�ZLR�����Q@�Hl\�{	;L���EQ`�M�mW5�6���E+t�A����1��X�
�4��dm6�#<%��I���e*��?d~`ͱ�;wq~�e����U������]ȫ�`5KZ��l �E$7>u��-�<�B�������B�rwiE�޵w�z� �M�DG��H,H��c��u�i-ƻy�ٲ'/��}�qeR�=5����y���o�V+P����z��і�X�h��5��/nRd"aZ�uF�t��K��T-��5�BAL�̲S(I`Q	�2�	"*Z\B���IJ�i�@i��t,�B�mʅE��ށ�0<�Wx�v�J�(0R3cdv��N�T�Q�WOo�γ�g�|�nt�䂴:��-;���ɮ>� T&}/�Kl*`a|lܲ���R�;��>��*k�?Ҋ8��pХש�ؿ-
=��A넿�q?�����܀&0��%�e�j.���, 	�Is�fO�o����1,߯]������H����t�ߡo�L�������bv�AՇ���l�6Eb#���5�! Y �n'��A�BeP�{����[�4>CYыL���!נ�Q�X�I��](��*ʓFҘ�RE��@@;-���-
���6��Qc�Z#�R֪�qT�i�+h�@�(�DBZnM��wߏ��~��ַ��b~~��9�sgϙ;M�%U	D�ʄ�X�r@A(!
�]Ȑ�X��b�f�5�=�i*�Y+rH��%-�Svj�����Z ٙD1���nZ�߅��T�S�<�/�����uL�R���L
%-�Jk�F��tm�i0%\��>�fǧ	DX�.���+߾O<s���������nʣ��?�o��!�w�cؿ�.��dV�Lu��r�ͭ��jB��D���)�ݻ���=��ԉ�8y�i�t&^ M�����C��G��m� 4�|� �d�bt��LsN���'Ѽ��s��5�'�m�]o����'�.�)����0��s��!�+^<w��s�J��[�E�n�
ڵD�D�}�Ɍa�,!N	��J!4>��g��{���cfZ�m�`��w��
����Z	��Goo�x�������)|�k?�W�r�!�y6�Bt�*�V��F���Y��Y�升^t��ڦ2+z��28�N�B��F���O���)P;�n��MW��Ķ�D=؉ D�{%.�����<�46�/��|��gI�u���ba6������������#D�dX
8��E���D���	��q�
��6���F�	��k`��<�����[���ͼ?�ə�z�$�0����K���Y�S�I�l�*O��Br�Z��4X?�p�N@�4"ey��PK��S[q��T!�2m:��{]�H���<�4�|u\��A���9m6ަ�;�A� c�K���)�y�S]_��	Sx07[$JˡJ! �փ�hx��;�F����9�dG]�	�(8ݍ2�J�2�T���
bb�����>�+��[�$1�*���߼�w_���"�a�KTK�KD��$�D{M��\�,�hP嶐}2������ZMs٤l�A�nH�r�i������h����<��R�ʆ<�g:J�'����9���2���p�|��Z��@�� ^
�;?�̊R��-�V�_�X��w��#�GUen5Em�emj[Å�S�����I�ރ
�ۢ����Pu�2�(_�Z7�mY_=�fj�*Mcݡ6�)X5.��0a�V@8ǖ]�a�@mz>�ˣWX�2�~7J�"׷\��	^)zY��֭�/��/�{�D�1Kka�����o @�����X�������#��Y|��sD�Z"���f�j�&�"�~\I�ͩ��Ț��d
�Qp�u!@��YI��}��@{]1����M֋�t�7���m�؀�:�D�<�π���*J%��z�H{�Ƣx�v�����e��.�����?�w�o�u|�/���=|O�p����ѧ�+��!~�w>�O��?��x~���pts�T*����/��O�Q=)-j��/��,K
�`�>ͩ�2$}hl�\�ܥl�ZS�|i�9�ҟڰT,�$�,�\��iYJ���~fXg�thځ��T)M���X��ZR�͆yB�W��$�&��K�	��[|&o���N�ˮ�|�eŷ��IŖ�R��Mᰀ�|�A|������|?�(����yTr4ݝnu�����7��$������ǟc#��jC����eS�~V�g�Q�1�Ŀckݤz�s�M��y�
�VGhSʠw� �-�����YZ ӓS�S�DI�$�u)ZQ��Ʉ3Y\���K�8M��@�I�M����w�mA����+���(S�-�fǵ2�����E�^���.�� ���hU��ߩ�����O��'���cǉ�Ȩ���v���$M��.)�T�M?�_�(�T&AX��ڶ|X�emvU�i{�xkk=�:��t��R�!�F��ug}�S:f;�adA��mDr_�Q�*Apӂ4U��s�O�J4��f/J%���2������6:�[��ϗ�MA%5��R��@��|�8�|g�F���Ɨ��-<���"��.+��B,���U>J"nAR�Q=�Y�/��SqGYI��[E��j90IW�`�h���[�
�
�ˊ���vb���>�n�ėr�5�͵�w��6gI��sW�IkS9�KP��O�7	7Y~|7��8�x��L��/����g��O_B�F�����P�9��(;T��A��f�=�ĺ��q��A�����sZuC��
�W��ha�R�
x(h��4l��ꡕ%E�%`TV��6ѐ@��ZZ9��o�Un��v�ܹ�bʒE��?��%�^�n��3I�����o#�SJy�J�Ț���S^^�ɗN�Ѵ}�&�'ݱ>�~�%*O��Rt���E����&�:sS3<�1v��k�f��P∆��=A���"�W#��<@>'��;ԁ9��\���%��|Q�"<�"O|xvdc��u��sXgE}����e�G�D��7R<�7�e�,�w�T�I�^*�֜8�9�W�%Ѣ��r��n5�G��M
I��}dщ��~����ph�y�ܚ�9y�Zo����qjꢂ8R���!�z��Zej�Zl�]u����wmmn:91�����o�����CO��K�S��ɖ���|���������~E6��5��u��狩,_$W%���J�m��_:r�߼�JjmuP]��O��YIY1Jr,�-%"w�b��H�D��8�MSoq�SI �b�(Eyk�4:��9ֳ$k@��Ib��S��A*ͮd�R u��wE��FO�� -`�t0�c���	:���d�3��n
�.]��g��O��Y9z���4�U��`h��(��:����6/��kеa2�᢮!3+��rs����-�q�}}��Մ������/�٨�.)?�'s�Vb�.��F��J�iY�����f�,��Vwݥ��^�-���Y.S��T���\%��״ɅF�G�(��l(1t�}Y��K��Ǝ=7҂�U�}�Ē=��Ǐ�/��_�����M�O2��{��5�Pa�kM2�I�P���5�Ht�,���Srb4����j[Yp�Ĝ��4i�KKҙO$���ړ�bS�P�VSW��ш�\%%�g�ϕS)Z4@$
,-S$� U�.� ^�����s�(�?A��7/i��׆'�X*�w͹�͏=z����Ĺs�
��1e��23Tv�N�(Q��?�FA� �(y������'~	w�靴;�-�ٞ��5�+����k�}����wRP���2�ܗ(�@|��
�0�Ei+U��/��u�V|�>�O����
vrrҢ2{�1:t�K��P�p3�J 3�Q-�x��\R�`�$Z��v^g��iwSx�̠�hY*�`��g{z��c� yIK�!@��*1*�ߟ±�g��I�k�A
M�K� ��0C ����D�ss���|�#/���.T@�T|E�@��V��/ڃ:eʒ�b���6X�*�p��]��ѲA�r]n�icY�*b���1��Awo��)�Y4)E�c8ce��蜊E�h�6e�f5�-�ֽ��GU{��-�����dm��QR�!��<�0�����fC+����"P���p����/�k%9$��r�l6���'�<��ZM�]��줍�(�>۩���n�q;~�ߋw��-x�k�ĭ�܈�o�{�݅kvl�����Z�u�md� �f3l�܊llM��h1Xe������Sy����DR��&LՂ��tLc�e�X���j��**�8BAd���
{��`C�>[k�i \�fa~��i�q�P�\�rW
��;ѿ��<DTr��,!tv�e�5�$�Q6�p��*$CQ�XtZ�06o^�[n������`��V� ��g�t�V���#���ބ�3Yj����$�T%rΙ��#�vV^+Vc�D��*�oU~֒�uU+.s��W{kgCy}BG$�2A(׮�%���țzM�l}�M��O�Ef�9��/���. �V+��3dљgO]@{����^n�6Ym
�pGH.Z��V��%��@�Ovz�v� )p-�$<�k��P�e�d��(44L��*��M�H9K�822��[�X�������;Ʀ��dIh3iLO��K���e�pwV?��9V�'����[���~�O�ɮ3zsP�!av��AdZ�T����h�m�T̂ӳY9cDx�q97�e�'���'>0�dep���`5^97������>�o~�~Z]U*�>ҕ��4ץ;H��G��i#l�:����tS��)�LO���NⅣ'�a�ϔ�Nc�����T��R@��`W��P����,u�?�|^���o���D�y��ƹ	��˗/�؞ܓ�O��3�<��g�Z��N�>���Q��tL�Ft������
L�dA�"��u�#_�����"K��e]T�N��γ�45��Q6�e��\����i�mk�k�f��<	K8D�5Ia�&��/��OP��4��MP(�ߍ��(��*2Z�����k�O�u�:xU*k��B�6�N#` @J�N�q�́���8��Zk׭Z5������22��ǎm��-�N� ��Ֆ�M�Z4��u����2IRǥp�;��/z�]þU��S�1@@!�nW��y�@�'���נo`��7������1���K��p}LA+Rx)*���1�Y���Y�F�7a9��KDAm�+����?��_Ǟ�ֲ �T��վ�H�۷`��زeV���:�+�VY���g���a�����$�	�y��ع{�T�l�}�,����ɏ��t�U-�*��LrSxj�)����jZvCY:��Dہ �)TXo�E'��N���4�[�c6%!�"N�7�A�.�'��MfUȽ&47�UˬP���7��g+��]���5���ig"&���T���B��:3kS>4p���t��\64�9=%r��J�?3�Ӆ�s36�r'fY�YwDl�v��$��/nlgc[����( �����*K�����ٮ��e��՛�j���֧m��)�v�`W�L�D�����Kh'�R9�ZՠI ��&Jm�@%��O�2@��-	��g	#ML��NRt��1TOe����6Y/v"у�b�T�U>����r����%
�dN'R`G֏��ͱ#
(���-�#��礐�TM�j��bcmT�R��q�m�]���?�[P	���(���	�j�Iϒ`�e�gJ跔eK(Ha��V��d~�1}.�q�Si�t�Qv,����BvT�UW�����_�ڏ���!��#�QHR�eL\�-��:�¶r������5:?3C��,&�U��hD@�H���Uڪ��$�3��xEOQʟ���	��U�G�lbfz�|7��d�
m̔�����P ��$<��s����o�N�ݩβ /\���/Z�)��R���|4N��d�S���jb&e�JV0GA�\�GqTS��]����Պ\& �"�\:%�ֵ�Dm��
;&m���i�6�@9�1-��?��a�N.Rv����y~���6A�/���J��xBnU�QiN��D�=��0h�@_�z�r@�,Z�@���JȪ(�ue1�@�{�m��[�y-^s�n<���8�,�+�D����Ѧ�L�`kS[��Z�5�e��p��������џ�^�z�����G˗����ݎ��j,�`{n���a1���	Ԕ5L` ��7R�H�����+���cϜ�|a	�x�� ��/�E��,���r��w�x�[-�}���♙y*�4R�y�93�i��~Z���

�BA?V�\�SgG09��W��ÎR��&�+���[فB�0��5�Q�i���Wm���4��URb�-��R�%�)bj����y��]s�$u��Vk}i>V��֯�����):L�O+4j�����#d��eX����B�ޭWF���nt���p=]�DJ�كd"���.
��1�惝�8�6�c��,`��-+t�0����4a�D�~��z-ɄEo���Xy�k0t��H�B�-�(h�&��Wڟ����>���6f���M@���Ӳz��|�6 -��f�X�����M$����-j}竬
�D뷛
�ZH�+�!��ġ�&t��(��m���D�
��C� 
�B��Sx�6��#��� )x���bqZ��J΄�-6��=��A�b	�1)��Q+����sXX������1�>���,��,H�SЈ���M���
�ge$$����g���>P�9��&$�Z�d	�M�:i�(�W�eTYg���'��=%�x	Ek�L	|o�WF�M	~寵~�{(8l<�u���z�kI�B�Ka����c��O����m>;_b �p��ن�%*��~���'֧����
P8yY�v�բ��n��Y��ܫ��)ѬP�,/�Vі�s�Q���5KX*,`��!Z�i��i\>{#��`���yހ���>��,f�gM�+穬�}�C�ȯ�
6oي7��M��;p�M�`xx؂4}As�ZBZ �A��EiѬF����dS�`�����t�I�-�SEޒQ�	�o����M7�쩙���E��XK�(�
T��	~��ތ�g�{��{��I�^a{+|;�E��8�i�_t�X�GI6h�xyΤ-�����:�n*M���zxN�ż|F<#���86��e٣�����O��u�:�|��y*�3�1��ɵ�d�Eѡ�"*5&'~�&���߂��ۓ�'� ��S�FߕGVcqz�x+J����|.mu	},9ĢIt���k�C,މs��8pb�������Zxq/e��~�ܫ8��O�?��B;n2���ljz������~��q}�Yd���~����������c�=�G}����=7�@�Q׬�C�v1]�󇎙�-�"F+R�~e������c4��Hbxǥ)k��&"��U�5/��@v�2���X��i�ʓ%�l��}��˻hQ['+?;��<�ͫ�)P
���1��u%�5oł�iN	�g�H�,C�X���r�PIQi��Y���Qc����f)���0=�!��m\*��`|j�sX���+rW~K9j�s��9���Q�wb�v���M�r�]D�$v��)5і�W�l���O��ZW
O��,��et!lTx�s�+���^c��fg���R�*���]o�}]*/7�>�-��d��-.eN/C�"�ǒ�"�V/���a��L��rF�+�<B~7"A7��Y�5�Z�Pӂ�����o��%�V�� Y乳p��Q*�"������� D*k����Nїr/ɭ�fs:I�꺎m.�@]�,�
�@�Y��B�EwjӫszJ��w	7>Ls�$P$����@������"!.Dl�Y#�,V��<��ma�z��4�$�HJ�_�!��g?����L�mL Un��su�놗�5�a��Ү佢 �̢ͷU��2�x�L�OQ���V��W^Ge�Q�x�as��H���_�La��I�)w2�WP�ϡ��Pwj^�G�}�-�\"T`������$A��6R��7���i;���/Ѫ<������������}�{�i�&;v���l���[�l�Ν�ɯM���%�߭�b��[�����$Z�̶�˭V��K����k�
D
�'ES�^�a5�ZH�X(������k�����xy���t����5M��Q��-m㜬��Ft����qk|?iXQ���Ji���j��-[�.M���i䱈&fKY�XДh�4c���R�f��/ �0���8�۽�a�|���K��z�-W��,�&�'^г[�����._gTi�;���x����9�y-/��Xd+<ڳ\���Ŏ��,���b�
o�V��&��}�$}�5=T�wY�T8�iy��(��ň�%(j��E�}fN���|�/Ѡ��\&��x䑧-븄��{WG���R�%ލFC|��!i,�KV�9���*���D�˛���&G}!�$����GA`a�<)�N�jډL��0:������^�B��VQQx��&S�!W-�wsY������D�~O>w��ő���xi� �3	*�2A��Ok���W1:��c����e��6=7gkpͧ�T�(?_���NKS��Sy
���6]�M���pST�Jڬ�)"U�
�Q����E_��/���(����P�՛��ŭ���v��+7���ۮ����/�"7� ��G>�u�����9�Yr���<me
�"::#� ?/p_$sRHԲ�DpV�Pw��hM�� �&Ok���B��iZ.�L��9�B	��ـ`� Rlc�X���O����;�{O>y��h�;���XV7���8R��ϫ�WZ_j���9����?Ȝ�Pk�1)3��I	
;��av����J�I(K�˅)7����5��ܪlD)C��ڕ���Eǖ�D7R攎<�FZ���`�0��q<��!����o����HWxe$/�Z�J�H�]bK,;V!ˎ�FП��נE��>�>+�" ����*Sy5�!�	z��GQ���*��fC���mx�o��uC��)�)��Z��/��o��փ���V&�o.e��"�4Ug�|4r�2�=����o����������G?�Q��g��������@��"7����E۲e֬YA^�`|�"ۋ�'؆��(����{�F	hSq���Td*�~�q�����sZ9*e��*-��I�.��N�,+��#m��:G����Ra�.<���2�cԋ���_`�I�I�+��I�S+�Q�/���i�ݢ���d�$iS3�kE*Z�嫟r[÷K��@&�w��J�A����2"�XHk��]�V�c���#/
�Euw��Ɨy�V"�$��**���p� �����P������_�]CB��?�pA�%�D��C�bs�<��O�!��!��y�c灤5���\-<��A-aAn'��r�5��X�{���·��ji�X� �����B��Ztt��E׃
����V]��t���M��7�zv��ij�7ծ	Lg�p���M2_sѥ��]�>�v�ue��/��B93Kd����[�ĺ�nB�oM"b��X�b��BM
��4Q�|����W
�NO���+����?��c�0����FǪ��bf~	������\Y��@�P
3��e��m��b�^P~P�4M��D!۷nv��F�l،�l	S<�Ǭ�e��8��aG�ª�U[�]���U���v�f��m���U��C�t����nq6�ǹ�EЭMϷqN�eE����d`� bQu;��L����U&�j�^V�]]a��JT�RdY�5GeWB�]%�
P Q0���nZ@d�\��Y�e�._��2.Oͣ��A��ë��+9�"1i}(��܆?��������'��i����d��=H��m̑�A
P�O���v�m@�ȟ�DMdm�]ߥ�Č<`�ܮf~��������K�J�wm��0�0o���
GT�<s��b)��]�d��x��۟�o����w��Y�/eJ)���%*)��@�Ц=G�VK� L�]Tvk�:g;�@ګ\�vC딯��M���7M[҂������*�RS���-�V���l�_������|����k�4-D*J>7����N��
� X�$�G���?���_��l�aoO:���eM\<��w����
���'q��ah�cjas33Tj�ؾc+��f�z6�������������}������b�Oc|�����X(��'����>��Ck��֗��F��e��v����&k���֩s�x��{�Ɔ5��ve)�S1�Q�i2{D�i2�?'�MM>�FG����l N��^"� �ښ|l�f�@��H�o�5Nlk7��VAՉRՒQ���e[�U(ū<dѰ�]qt�x)�Y^)8љ)�]P^S��:A�)�"7�ޥO��"��|{5��͙N�{I�F�d`p���+V�6�i���ݖ6NSUd��Gh�O��k�r���2e�9�&!��vZ��'h�>r��Psd�tq���tJd
����ʹP��)���p�	�%��R�]�7��J��&m���ШB�t���ٜzi{��r������uN��V��K�ІL���R�%*~B�kw]�����P#j��R�U��Κ^Z�MC�*���)8t�^���3���h
�.��Թ1���t:i��>�#e+kXa���]�Ok�EPUY�*C��Y.�5���u�y:֯�\��E��&�	.���[�L��Qt�Η�.]�S�r��-�b�r�3e�	�Ke
�)�L@@�Ջ���V.���"��MQ�*����{Ȥ`T�^
/�rgQ�0��r5OQB$D��:�£������\�Y̡H`��F��Z�	�4���E��淄��l���_���g��<��������-�����������w?-V�TɅ��_�lR8��eu���	L��:���.���A[�����G!��!%ט�����'��Yxboޯ�h��Ss�4p��,~��G�>HZ�̦���e�6hDm�'O��x'��;��'Q�l`���A�Q>ǩ�h�X_;�����S���{
�w��=,�2~(�\��q�J�~�Z��B;��1��E�r�"�A,�fٖ9�mZeZKyXi��Nm)��ѣG�-sZ�f	\(�I�{��J��o�U�;��,צ��rB%Z���WBx*�j�@z�ඛwӲb=C^��э�+����/Ѥj��# 
Q��O=�2���e��U�9ҡ�?��>� �i���,��r+՗����p��wI�K��E��j��ɘ2:�}�
,�Ѡ`�t,H��vU���g�K�MA�g)�-ʵY��U*���,�VT�xREۣ�cǎ`zjڔ�֭��G^;�]gSH�����X,j���#��A�=[�]�;��ܭ�09@`%�H s|�
edڎ�Ư�W���5�����OO��tz����9T�]����Bf�N�����b>�BǺ��=�%�Q��&:(K}�P���r.]���q��*� ����"�sQ��3D%ܰk'��{zb����?�ܾ���!�`eĐN��u��@,�<rRI�1Uܗ�~�b�!��)�&;�̶J���:��Kǫ��?k\g�o&�����s��I
m�Mv���/�+d�0��=��01Ų���>�$�L�M�7�R�u\mz-���J�5���l:mQ��\��DK��6���DjM|�Q�_m X��Wa�G�؆<�G[�Jl���Xw�=����x��9��4n��r~��Ld�	�K�h�q5��ry9;�=0Ծ�{Q,��zW�T�dHp[+�:��w5��������U�K/�;$����*�JӠB�EV)dq��(;��5dS
�A�B��ƶԪ�� �+�tj�]ؽn��B.]�B�܍���хt���C)S�����|>����`�)�y9��.l�}�}!���5o����-&'�z��f�������Ocjv�d�-���ɣX%�s�-]�m�:J�/@+VP^m�����17\.c�}�RѨ����)*E�JaH�	�*�E�
 j&UE�
��T���e�o�:JM3e_i"DaP���������[��82E*�py8��\�\�e}bpG�h�u��'jv�����+![�)�Y�GJ�L!:��"��=l�\�}� �O�07=���Y�c�ه�%��rƵ�x���7v!�zha(�|�q�9D�x]�t>������,\9m�؏7��X�z-n��&�u�ص�Z[a�������k��7���r��ؼ����M7݈m۶c�ʕ6>�1L�A	2�=F�p������}�b���jF���w�鉀8�IPVǊ�H��ar�����B��H7�硥�C%�`;L#M�z7\�[7�0Ӱ�ً#|�YҦ� ��Ŷ[�P"�UDy,F&5O�<mK�-T���2C6O���.R)�Cs��uи�ףu&��t�x��yJ�
 ���/�*�%��VD�E������x-N?���N��4R"����T��X��|�h�2�P�,�ߔ�<Je��0�$�%O��y#����R`����E�{lS�y��q>�����26��N*�"�-c�M7!�7���9��<�s�3��qƇ�� ���W��(������{�?��⑽'ɨ[ V^`ǰ9�H�j9���X�NZ�z �bg.N����d%�t�8_�Q��w�?��;,��I����0:O��+E�L��b Ei��}�6D��ZN�`$����r�1,YA��V��4�,G�y(Xj��vm���Y�${}q�PĘ°q2K�JMs�zz{��;`�*5����(�x߯�(l��L�E"�ȴWG6�"Y��t����Α��"�Y�Nuq�8��%�U�%��z��ڲ;�z:�^�2m�헣rz�	�|��U�Y��~Jy^݂���oG��J�\
�OA)�Z)�̬�ƙ�jk�N���ݜw��|��TFe�$�^���g.S8;
I)��� �,Q`��H�Ά��S5����k�b��A�i��(JdH�i+�G�mTR�)'�[XW!����_�>[�4�����=��%p��%�lZPs�r�*��
��w���4�l#~>��
���ݲ�3Y�G�w��!�zT�7mlEA)�6"�L��l'ݗ!H�bs���D�N�"Yi�F�/�xӼJ�������������o>���c㋼'I�A� "G:ҧ+���O���h�\�]����P��",�ZӅ��V0_�+���%㦀U0
�Y���'��y����B돂�nB9�`_��ƃ.
���^ܲs�"J��$ܗ.i�V
�R�VY~�g�b�*� �M�k���?�sX�r�e`Y�j��~��ؼe��/i�2Yw�r����w�:
@Z&
 ���6�G^�����9sSS���2n��f$bI�7� �p�
���_ -��im����a���!n���� ?G�!p_%�O�L��� Ϳ��0<L�I�P�9x���j��-s��[�D�NJ,���h�#�ə���:۰L@�9�mm��$�Ri)
]92٩�7�Fe$Ӑ!ɐ��P����J��꟢{�b�:V�u�w��k6��3T2S8|�<��,e����hO�}f�e����+��M���!%!�ۮU��n�e��\<Pd�j\��	�/XEI'���$` ��+�!�x����cG����UĮ�ǚk��J�������jW;��D��*��
:b̄$w痉��M'X�r=��>{�ز}�ԡ	{!���ň��$���Og����U<�����44h.Ũ0m�-8�;�M��Ϋ����غz��k����b����X���Y��4�&H���G��5X�}BCkP �)$�HV�>�ͽ��J)W'[^CvRS�K�D�V�r����@��@�h�)�A��9%��;J˒V��`�H`��`��߆�ބJ$��<2d�W��[֜�}c��'��>��~jӍ�v��}��ܬ\z���[�B�r��d��&"D�^"A6,��"n ��
�IϣZ���m��G��i�O���2si��im�E�D� i��+f
2�"%�]�Fɨ���6W��Yd��
ɰ��,K�L�䏢����S���w�v�F�h"S���ƿ|������2�����g�?��T������C�H6�j(���e��s�Y~j"��/�@TVEc(1�\̲�ñ�M�ռ5�r� ��+��B%���Ij�_��s���\=z��BE���}����83��B[��#��,���;L0E�����V�˛��٧�zZ�MyÃvZ�J	�%H��{�^̦�(T�'�����0x>E�15�F���f���_�&�˝��/ʢ��i��ǥ`��� �Ǉ��Pp��(���\��fgg,�r������߿cW���062���	
����k]���*M'��YҖ\�gN�ǣ�>�wy�������<�,��� *�96:��������j'fSX̓wI+�h�e�i�m5߰ƺ,��ۡ��S�D;{��'�./R�Ϟ#8QV�ܶܒ�jni�
M;/�i�S��ݔI}�z)�"(��̢���y�@1�o�הr��&M��G�WZ}>F��C�уvOLkY.�����e�P����(�z�b�u��IZ2���
���9��$���ٳ]=i�G{}�C��*`1�ri6�����L�䰰�U)<�j0]�+��V�Ob��:�d��t��"}4�8�i\���21Fy<�b=�@>CP�g����T���ӦiJ�e.�{?y��yZx=uي�Y-�ӆ��I�c�i�
�LON��*��\i	'Ό���`�X4/i�PH`><��38x訍{)Sᯡ�F��ڬ��;��� �(T
T��Yxڭ�/�t��kVы^�*�&�EH{Y�-���9�Mz[�
QkB�^�I�B�*&/	B��2"��W�%vb��I&��� ��k�
�$Hǚ˧�Bt�fP���+���Z7,O[� ������v���kn��;ތ��{P�v��B	���<� �����ML�Mmg��6�O��ygo����9��jg�.��tR�g��&%iϵ����J��Ԧ�t�ިb���f��h��;�A���đSlK�8�A!�n7�0�GQ��mIn�ȱ����*��Ut����T�*-A�t/U�;H��E)*=�:Wn�X*�OJ^B~l7�'o�� !�JaͤG"�%* �d��I�~?r�� �G�v��K���8�$NRp���!�<y�Ɗ��@:M+4����<���+SHUXI�5�@�%�iUNC��K�_�V��ɸ�d��-��!�.d�8wi{�?�'��}>�o��A|����عK��{�\a�&���8ru*wВ=��ȽTFKT�K��dɊ?-�<i��s��=l��%�4�OZVa
\���XQh6��m��h���+��<��� ��GsV���&�Tyb������Zx�ע3B��!������g�GGW2�Y�t�N���N�8i�{&�z|X�z����'l��B>�i���1<�)rP�R��[��ىx,FŘ���5y�۸yz��p��	�Ѫ��[�b�I�E^����01W% [EE���	�kP4�_	����� ��yO�^��n�~V%MONg𓇟���"��NZI��ȴ�4H9���0����ͬqT��N`�$�"k��W�K�<��&�D�!y�<Cep�O�
�"�hӽf-��I{�o��r�.��`wv_��<x�q�K0�!Pk�Y9�M�o'ЗlW���3Ey�H�Py*py�Vmפqvɲ$�h���b9���@Ph��(���T����h��x�-2�'�*2S+�Gh�%	�z���=�c�|����$�\"�vњ�K3�!�H��1K&|u��Q0VP��>�粖&���3x��a��.��'�!5RBL�cY�G���珐1�:e��b*M�5��5y|;5Ƃե�x\�4$+��
�E���
O��\����U��\�Rz�&ƚ��oY��B�Z.������i���^cUY�:�Q�u�+�¶��6��r�BQ%/�Vx�P��Le��F��#8�ۯŚ��D������4Q�)!Ua\�Q*-��X0U���N������Y��7^���\��F�OB7���5V$C��z�>[��4ݫo/��N_��ri�=ٓ�>;r%2Kgg�2�pv�L��|gM0ʡ��6N�������.b��!�Ka6�G89H�b;Ө�)��B)=�o���^>C=���f�@�@ڤ2$6&ck�����HD)�F�<�>d��HlM
�&�[��j!�(�G	�C�������\���Sx����3q���x�
�g�ɜ�����ٟZ�F+^���gi!R`Hi�������N0���.���ǟţO��S�0��c��7~�����S���TR�J�H�J�\o�'���*5��H��.�f����
�C3�\J���Ci��vn��f[��,+��V���JC�i'8(e4d(&��;J RlZ����-�,Q)dQ�ip�RP�;�ʳT���v�: %�*G��O>�'�zΦa,�Ob��>�h�?v�9Y?�(Ju``�&�/,��x��Ec���d��F��N@���*C!�2k�V*��>�};�޻�l��p=V�4/���~�(��˴�f����.��Q
X(
B֝�C�W) %xך�!^׬."�8��Y��kI���x
�>�4��i0J������KY�RU��K��(R^���+�^ �ҕmG�]"ߐwd�ʫ�V*;��&ϱO�� A>^n�T�y.Ҿ�`���wD�ضi�l*u�ǟ;���H�@�O�G��w�i�:�{4�*oI�e���5�]@Gr��!��v�<�f��*۵�4�DF�KI�y�%��P�֩{���z����,>�/���,�1��P�]�TZ1tQ�H��<�-�|s)��y�r���o����v D@q��6��f�9O�ns���W�1�6�S�!
���
9"��{�l
�G��g$⦠&I���d5v/Q�"��2B1>�����J�׬���0@����s�#6����+��2<}y��Ke�juP������|GT����"m�o"VS�%ԥ %�}D?R���\�A֩ǻ�Bz��y�3d���3c��`����(��kh���S��C*%cH(�4���߹F��Y�
��|.[�[V�ڄ�SQZ{H3�,:��8�"|y=5�����/��Og��i_m>o�0 �%�,U���lVd~��lS�ؿ��^��Λ%L��]+H�\�K4Z+�G߾��Y\O�s��L�^$�&Rh�BqhjM��"&˗���%��)�O G�����fpt�Ûn�@��'���_d�ݖ �12%�eg{�p��	��w�H�ʄ
��җLRHհn�L^��X\�i1ڀ�<JcF�L!ަ�=
rB����E!�.��E�J�B^���@},~Ҫ��h�NMZ���Ҁ�t� @�5oI�o�����S�F��G(Z).*`	� ���Qtb�e��
-Y�\��(�A֍V���ĳ�HH�U��yJ&
%��8�.t&��3��Da���&�ݫH��X$�Mtк�\�r��
�H���[�&��O��Å����y��/�`�ʢ���sW�T=7��]ߍ���k���K1߰@�{?��Thac��$۳��p��刍����{03=��+�L����ՒRe��ϱ݊P�Pe��q�8!`�6�"��ڽg7���q���i���/^��_��_��u���0��S�{ ��'��հɴ
ծ����Q̚�(�Y�9��𢚛E9u��\�g~�W�3o�պ�ҕ9������-�B�~�T.*(%�`�TҘ���S�.!#H�:g�X�Z�
~� ����I�H�-5�Y��]�&���ya��0�M*/ڔ���!����s�x߻ߊ��O?osk�!�7_�T��9�E���1��<k,Y.�BJ���cH~�ƪ��F�2aҲ�ݑW$o�-%,��$'D��)���R{ʛ�f}V����	¤�S3�ᶛq�k�����������b���cC���;0�������{i������Ә�/!.�2_:�QLRi�E�k�����'���c�$e.� @�Z��+�7��ef�(#4�F#טX4ց�t��m�C�(�fL���>!jE	E��$ղ��6	����O�Z�ձ��Q��)[zD�<^c����M�\>e�mw��W�=�[�z遨��c^�#�Y"�t�"��o���\���Zt�ތ�5[h��Bt�F��lFr�$�nA��رC;�C�����X��af)���)����X7M�hYG.S�B+��""omv���zs������S�9J�_�˕�9Bң����qW���lg��lm��I���W�tN��R)(���D��p��YS��7��l��Y����1�<�r�]�����mQb�;xz�R^��V�E�
dz�BZAʂAa,7�V���Jb㪕�En~Q	j�S���l�:�۽Y�~f��Ac=hI��yi��q��Ÿ�����3s�b���(]ާ�g�Q�{%��k-����K��]���<&�3����UlM��J209�&?e��J��.Ur;���k��� �@ׄ���4V�r���7�]�#�V�T�[�@�b�2�*�ZH�D~��U������ذ�nZg�W��R�\u'��X�><�@"����S��b>��$:����刮�0Е����fj.���Ba��k������q��5���z)(�dI���{.LS�Ż��fQ� V�\i�r��[�\���=�1���Y�9}�ʌ�:1a�#h�x �󚷥�!-J����{n��MY>�&g�̾�2�p-�pT��()�^\���OQ�����2����5TN�df��^X���ů`�r�
1JC���f�禱T^�[^svm�q��,��IK���p_�i*�f��g��iv��?��h=I7�A*��2��9Z�T�m�Oz0��E_'�q~�+GM����9���}�V�u�x	Ȫ{Z�Q"f+����Nt�\�W1ܟ��^'vn݂��?�%��!�Q�"�qv)麈��(���JE����V�J��r;Q�&yLi5eD9_C��]�4UB^�#SI���AFA;�~
'/�B�8�������q3V�YIKϏ�#38tz�Y���`_��Z�0۪��k.�(���3��_~gg�0�a;b	�i�IX)�L9'-a'T�jᱲ�4��d��,� -M,�p�<�Q��v�ɐ�Ñ$b1Yxe����0�&��7�X �²���
�u6	�e����xU	���}y�A��|SQ�S�\�X|��S���v�/���ޭl Mkԧ�-u+yv���N�ؠy-w�,B%��3Pʩ��R�x�bO+�ƅ�i��
��������S
SM�������4�"Ed�/��`GXݔ���ݕ��^� *��̩q)[C<Bbc�g)\O��s^��.����ZϓPkm*��^��*�B����T�<��� B���[n��C�����,[4�-D�qS`ש��lX	oi���mNPL���Y���j�æ]7�����Q����"���&��}�o؀ͫW��ާp��)jȧ�I�cJ\��7�'������ڎ�m��C4�(3�C3�H�`��%f�@��$%r�Q���Y.-�T4�V iB��³g�|�\Dr��qe/j�
��H=��Fe�JX��і��
�T�lW��LC	4UXY,��1v�
D�-V��=}|�&лq��{0?=���VK�8���ڈ��S{��Az_�C�}�%�J�ۂ��TY��t`�?��>7����8�;l�\���K%0��k~��E�j�Z��w���s��翏{��|�~�4#�2i�NΞ;Ks�B�Т܍ra*�z�Z+"(ף�l6����`�^{�L����g������a�&��.�����K���~�?���M�����'��+���F�2 �.b��!D�U��;���#BK�{pf����C%=�S�����h�G����|�ݯ%��m��+�2�tg��K#��˸Bk�Ll�-X�ZK���.�ْ�{v.e�w����j���,�����/�f 2���>�t�֮n��	ǅ\%���kV�# ��l��TP�p�/]F��l��OKPn�ɩY�*��M�J&:�G͒��Q7Y��~��2h=lMᚙ�f��F{�;YgZ���������qmS�^L��Ƨ�6^	���4vQ��{��n��!�{�4���c8>B>Dp͖.|엯Cw{����ܫ���2�{�"`��Q7���Y
l*	GZjL�e
E��V�U�Ⱦ��J�`�\�V��Y�02��Q�/R�m��㚭l("`�'!�dџ��-!�lR8d}			VԱ�(��� �<�Kcofͼ���_��~�J�R,�X"e%�����]��OH����D�0BPp���kPNkݩ,�v��;g�R�L����T$ؾ�:ɑVs�m�(V2���nB�U0�-����_�����;�ר^��E����h�R������j:��r�Z��"^�=I9����T�����L!��8�öwۘ%/ۺ��J�|��\�-��t�� ��@����179fkJA�B����=^��*���9Z!Ңn��E� a2��e"'��2P&�dpw�:���N��qb��O��yeէ����yYzdZ�r�,	<���U��&�:y��HK*Ҫ��Y��kS� ܗxL�[��0ܡ��O�AE����,>�Ϫ����.Z��w�]ёRx��vt�[�z%��YZ3<FRЅ2����7]ݽ�R�LLM�"�����v|QҺz:i9�0r��jKҰƗk�>��:�m�����- *T�f��`dS��2��R(gX*���)�K}N�����ȑ3��ݸ��6�ix��4����(�\�	��T
��أTm%ZUJ5�2�C�N�PT�A�ɓ�1ze�2Lc�M$�IQ!uR�*3���N=�L:��|w����4�.G���ѧ�Yd��u�����y�n��;�(|�Z1�C<с*�+�ll��/����5X��˦����E���I:d��V�H`ݚn�f��*�_�!'#A�FV�P'֭¶-��j���!$b~Z�n�Ѣ\�b��c�������V9-�K��~Z�C+��rE/zy?\g<�ޞ�4ͱ��=GP���"TP�q����U�ذ~5�r +��X�~���B���a�
�����>�_�
�W�5+p��-����c�V޿��[����&��U���T�3f��t%�b��=�����5�^�\Q2�6#E�8O��Px����"�ew?�g˭���bt6I��܈_�(�^(�P"��q���2H�2���n��&u��8I�dx�|�5�$��j A!�-Y�W�	F�z[�y��_'�����{���l�M�H;�X��q��SJB�<��,jw4ɣ�
iv������d+8(;E�o9	��W�����
C�zo�k��$)	BkR3�(��.�H����DwZo��ox�]]�&����Cw�<��B�����^�������|�K�j�T�,�2bȊVre���tt��D�y�%o���V��	k*�|y�V��<��b=�3�mȶ�-��zԢ�4�4�8O��:�UF��
�B�bhP�M/�pyr�:��?n�l�Y��,QQT\8}~�3D��2Be��>~��C`L��b�VD���]�o/�5�V S�e��:�<ʚ/��R�L�@]{�e�&��D3܍%��_�/�S��v�3ԃf���b�鹞(�ܵ h�M�1�*?���2���֭�'늆&���ǳӓ�FEX�H{�֤�*i���"�S5���avۊ��])����i����������<-0:���,@E*�%Ҿ��RQ�
ŗ{WY��R&(�%��[��V�и��M�	�q��i��G���#�����7�t��M���Hh�R�e�d��2TzR�SSSf�i��'N���ط?.^��a�'�T�r���>uL�F��TP�3��|G,�	�؀����v�B8}a�r�=+� _��8���h��J�(-�d�2j��´0��U`��Ƒ��y�R�%b��J-&�,�>�C�l�S,kH��5[��ʾfٮm��R�<F@&��qa�����ȏ$i�\@� 7����I%��ӏ�>*����(�-��_�Q����(E�~7���V��@Ѓ@ȋ��1���Y�n�I��0�ܤ�\��B�&��rO�P9��%cY�X��!۩�������u��r7��#C������˺_"�������~�^�L�ʶe"�%5���a)�m��I[�2B�vM Kڷ��ϖ�cY����񴢸lEE�5JEAO��5�4ɱ�YH�]���Z�����]��g:�y�>Z�\�*�"�d�e�-<Ei��e��a,��
��ė���m�-�U�ϱ2�?��~��I|4��s턑=�O�_�N"ZG���)L��.�S�	 �2���vT�3[ŗu1%���ٞ��U��C�z;�ea��<�r��-�Q�j�Ц>��rv=��sy�&/HB�P�1<Z��_���,mV�e�?�^jY�H�t�9���:�H��ID*���ѓ(/�mp[��zvQ�H�k~��A&��\E������]�6�H�h��+B�zv:ǟ*N
ZF��ܰ*����)�� E��*S��-��$hh1��E�֢¹B-��&RSPS;X?�[�4�	+Y�m��o��7M^���.�!��<��~����&�/�Z��K�%K��u�� �֚�r56�����c�U*`y�YQ�0��(X.�(���%T�k� �T�BH/Z$��2k��륕\�P@Rhj~]�t�����~7�2�i�Њ�cc�iE��s~
/�N��"��Y �U��\j��&o"|.� �"����Q΢7َ���BwT+���Xv���������JMQ���fh�uh����V5�p�"�SF<��i���M�K.�ܻ� ��2��Q�]�[�ߍݍ7��JZ�	Z|0-.�	��۔�;��]��H��|���H�5d�M����b:�r�J��Z���,T���h�Sk�K����,�V��N�?9_��b#S|�������Ry.a6[�L�dnǉ�(�T6�J��y�>?���T��#o��
����b#��g����zm��v�*rj���{�J��V�.���f	:���������]�UXH�!eҽ<Z'���+��YW��)�r�'���|�ǳ�xe]��H'A�T��H��\�#��>��Д/�O@�#��窬{���U���V�P����IA}Z���������^��E����#����u몠-5_X*�}86�ß�A<6����&\�
��Iin�/�\*;�,Y�ʨ��jI��i��O���e
N2=�)���9�'�KF���$�ga��>��|��?��ÖI�-�Ǥ�^����.eq�&�j�x��4M��X�0ˮ�]7�P9vu�ȑ I1��2%Q�%˖��8̳-�
ϴ�7�x���m�
�$+P)F� � �Adt�����]�n������{� =���էϹ'���{���R�N�jV�CD #�!$����F��L������Y��F�R�:tW|CIy"R����z�ς����f�^���\+/m��u�w ��J��R��P�����aa��gJ�M��{��~ir��D��)%�}+d�B�J�,�J44�t�W�9C�Jv�s��w%;j�+�{]*�� }�,�T�޲k��-�i��>�%��5����"�\C_��]���9Ұ/6Ii�-�J�R��EEuȤ\�"�M�0А�����=�L��$�<'�����`�a�Ԗ��ŴxA�U��I�EZ-y�̧�g���D���QD�l��W��S&rx���6jx\Z�|ʚy��<��۬YBZI8Ȓ���!�\!"��֜���h�Z}� ơAǲi*�4:��������ܹ�B��c�)`<x�{�Ѿ ���8/���k��Q�^7�.���l��CJ��:jL9Y�����JT�6uH��8*B6J�������{�-P���~<��g����Lyf�N�o��/ٝ7�(�����?��}�8<*徊Z����ϟ����a��s��_r��
�B1ocX��[��曮����a>i�V�Ο�h�z�q�:b�1�Ї>b����{N1\������O��G/Zb�z+u��Ar����G�ui(U�/<s���� �G�׶zmǦ��mr�`���\]Ố/��#�g��L;��(&X�n~u-�	51�l���o�7�Q���݁.R��8�56��ܱ�����{�267����1�bU��m��n��5����ɱ�/���U/���n�Ãi�};�G��\�n/u�/m/����w��t����ܛ�� ���o��vpUʿ���E�B�N�min���N;ݮo��X}Նml�"�����[�ڲ�}\�:���k���d�έ��;���OnZ:{��c��.���-��^���^^�ۿ���ٓ'xW��4_y�%�	��GxZ�) 묠�Z�G�u{e�/�Ր���\&���Vg1�����4&&�TV;��I����IxLm�h�$�;��/I� a��%O`1��v(�@�#�N��V�p{h�bt2�]x@ #��s2zC�B�UY�r(qx8.z����U��w��ߜ.���@�Q7��/�&��n���侅^�L�j�\�х���a���)��:#����M��SJ!��RrK0x�<��D�8 pivn ��A;�F5���p%�D�W�m���eqF��(�a6���y{���-���9�~���̚��A��C�<�Xa,�X��='�|z�h՚��0���:�%�=�Q	�"�B����ewk��]i(>�ֲ~��iKY��0����980�[.�M�Q�±]��æ��%)a����7\���S_h���������P�4O�9��f2h��]����ʺ�5څȳ,A�\і;�A��=,�!EO"R�U"J�Z�G�w]��J!,������P��Q� (-{�"�UDp���/��j^�֦�?�Y(�G	mY�	��Ե��U��yTPi׮5����jD'������O�c积�ISAR�G����m�7����-w�Ů=�h��|Ү����@����>H�7�b<�-��ga�M[��֚C���҄�A�hE��DFHx��}����e5������k���rv���#�3��q�/4�~���/n���I䮲�~�}��K��+�Ά��E��q?
�����p�5j����E��ڪ�G�%�S��	-�#�nC��1���R�@�e�K����^��MNL���k�߃DV ��\�VBpiG>r�'�s��b*T,r�JN>�K5�1�Vߵ��[���|>{(K�QT_h�GC�T��T����E��:�!`(m�W>%��Q^0U�NMh\����~������$||/C�Z���C�(^���U�J�?h/�\�c���m~�5���~�N��W��Pۧ�>!ɅN#SψZI#IC�p�����h+qO�����~�ڙ���Ԗ�x��E�� �9�~x���LS�Y�9�|���=p�-�`�r=�=����Q.:�*T/���>�AS�BߓY_��0���Qҵ�a���]��Cޙ<y�
�|�gݧ,
3Z�����4�=G��ς��)��������'^�Yv��5�8�� �b���?�{�Ր�Σ�H���еz�w��!���;�a^�x��`h:Q%`�����%��ol�����ت�mj�0/�C��ʮSv���ZS�Xl�A���b�i_c�����j)*�4��`٠yB�}��Z	ø�v-8M���m�򨛢�ȹ:L,�؄�h�;�*o �֭]لQ7-6�[��0�����v7,��A�(������haέ����u��6��-� � f�T>�K����u�h���W�2B��MO�l<O;+�v�Z[�h.�'c]ژ��q�;���֤.�ꦥ`�q�M�߶�b�2���`�ն0Lʖ Nqڮ����"t#к�A�sx��E
�;���x
>Pۀ˕��u�[F`�ch�@an��w���2��q���T�Ċe���@	xM�h���k����I�>��d�j����m��I�رv��E�ޭZC:	�V�	D
���be������>�qۿp �f҇�C�{��,�Y�)��jB�zT�F��vH�Z`�N�̷C�*�<����^��3��-�����fg��+����n�U��aa���r��Cw.FZ1/�Q4�F�fc��<����loY!�Nl|l�2�"V~��A&W	Y�q�qrr�n��Ʀl��²HW`�1�;51����l��_e�V(4���x�x|��"̡�#=��,�jk>���3ȍE��
ƒg�Xa�Zˏ]�e:o��$V�5������y�4�1���y��������O}��3��<z��(��hI�Q�	�8P-!+f#�@�q�?u���nV�����rS�x%i��ė��39�J��SM�));�S���M�
�V���5T*A����w��C[�(�b�7P�8�[�^�Q�Ƭ����I�t�F�(8���g_�Vt���䨆����P���u���+ a�����Wz#8sP����;�7�C�G�ŕ<u&Gu��&�8�pA]x���@���ȕ]�Ѩ��_��p��K���y�Lʒ�����K�X�rc� �AZ:x X�����V!���Iq������ʲ�@C�4^��m-M�emv��`o ���G+�#�ı�q���d�7�D��{]���"�\L��ڄ�Ѵ��:hUи�T��<����T�.w��v}��|�z`a�:a�i����p�N~-D�f�,�:<@h�)#����(�i`r`f�&�h�<�#t���I�M,>���1�B��t�v����X_��m�6�O�Ii7y����D!�5���C��O�X����$VY��&����D.÷�!�00���<J��Ofm� F������<0��ٱ�o���FW�hG��$o,;XH��C����vw������m�X� �rlnR>.W���	���V{w������5�U!�$`�	k5:۰F�
�W�1Y�a;|`	a>��B*+
Oʺ`���ƶ�\Z����V��/���O�{��%��Λ��%O��(��|�hm�I�B�i�x�F2�X��s�8gQ�4�ܴ��M���`M ���&Ju���֦�B��)����h�&kkE���#XV:c��۷�Ç
�,���Zީj;��M#0�^��P��Қ2�����Y�,�&u�Rϵ�mK�T*��lanޮ��ZˏYi}ۚUM�h� -Bk��# бq�#�Z�,<@�vyk�P�����lf� ��z-<�R�p�\{2?i3KW���a�'�c=nU:֋f�։X���&�@�8%�"�7��n�i��V�h�_V�β�<�4���,8��2#5/�aM��n	���V��\���~0�Q�@ےƦ��P�8�)��ɹ�����i��a�KWCI.���	o0���F�:\8��{zhs�A�	q�7�M�(�2�XQ��3ʏCC���| e4��ә�C�hJ=���O����nͪ`�ڇ�y��&�f��<#�Iɑ+�ß�:����([�izh�=����w��<T7գ=�����M����� � ���C�#ɰ�`��D�&�'�V5����$��3D�)<�N�� �te*
{�6:�P}C��Z���i9��h�m�Y����x���,�S4_�\�`]�e5�ϲ�5�F���uvf�;����jլ���!̼b1g�\
�ㆹsO!�4����b!�e(�"� � h��M4����w	i��d|r��\@�X�[@�r��β�0�5Sȧ����"��-���;Q�D����[�pW���j�-��ha�D}�De2ʽH�eYfh����	�*�)O��X����iH��P�$u�Ċ��a����0�6�,�G5^�{`�4���s��/ʎ c-8[���Z��k%	!���|���n�J0@���{Ҏ;n�����o=��x�F-";���8��`έ���;r�a���[������ہޗ�oCqK�	)���#��!{���d���{�,�Q4ڀ�9b��I[\Z�q���
�� �	����'�ƲX_c,!��h(���.�A<^��^\'�tXbs�����ɨ�`E��$��ߵӀ�kG-�Q�
���-�G��?lK�����I���r9��
��~��2����ժ�P�`꾈"��v�&���PaF۰�ʠa���z(��k���B��iOxE�y+��Y�KX$K݋K
V�w,>��f,!�~ɤlΦ�WvR�}d�G�2)iT��]�}��6ׄ8܊��h�T�֡Gk A4N|��+mm����*P����{Ґvvj j\V1��H�h-4�҆�РV���v���$T��>u�q^��
�;�,4!-$|�!C��n2��J%,	��:��LZi����Tʦ��?������:��<;���y��k�G.1:3�B����V�uZ>���G���X05���A�|X���Ԧ�b̂�H"J j!�
�#P� Z�#���;Y!�����H"0!툜�i���~T톗�3���G�A>qƨ�b3�(%fK=9B�ζ�X����`�I�y--Fhy;%�~�.�F�&���Q�R�yV�p��⹴��iM^B��m���{�o.C{��{�jXAm����k�B���X.�`'r�mK�CS�i�\�+�I�
ӇYAu(C�"�.B�F�!�#9#Sp[s!` 
b��HZ�'�����_�ȅ4zo&x���:�F��K$\;�jMkʚ�'�w)���мVM]GNN�H~͉��Aθ�j�#��(W���SC~�4��}ٺ�E(G������l��^�R�&%�5Ϯi�(��úmc	v{u���.�����F�)��`����עm���!�P P_��Cam6V�A?���ǭZ���\!��0����E�R�5�� )�M����$�p���q�O!��-
-�	��䟰S.��Ɩ���Q{��1��"�%a�����I�ݱ����z+N�����z����	��BZML]x������{��i���*���rK�_#?9=���\�t�o)�j�s/�_~��a�W-$I'��Č�O�UNN��+�x��Vo���Փ������C�^iч����P�^S�14wCC;�hx�U�b� ap��CBEC���jh�.�d�*MxH+�م�4�U�W�WM�I�>R,eU'Vq�)�#�EC���Z{y��C_5p-��� <��v���9��E�mO�d
�:_�ޱtq�B�g���VT����h8ɻ��q�wއ�w��7�B�B���{v�m�Y�,AB��[}p��wj2Ҁ�&�i�Hq���y�g��FD��S�#��+��iiCKm{����z��f�-N�kX�˫3�B��T���ļe�����S���wW��@��,E-�n��"�n�����|���i�1,߈X�U�}��y���ٍ�������M�k����P�%��IK�rO�5�JC��&�uH3͠^�~}�f�q5�5���k�)�	y�����Ch�h���0Yq�bi�@�q���I{�ՒC�d�i��F����謈-��e���1�a6
«�:)�E�F ��[\�a4��"��I�Ü%[郲d$D�PEm��0���)�!/ʧ��FVۡ���k),:L���EZ!˄:b�t���Ί.b0N�Y*��bj��}ڒ'�(��l�
?���8�W
�F�h��Q>����m���l[��U�7�I)@�	_��AJ h굺�@�^S���fƝ���K�s�&��̣��#q�CA4����a;�Q���h��.@y�./�jK1	�:29,�ÌA�p/L�
��JQO�i�]�8�Ǡh<_�Bѐ��NM8���4#f$�w��w)CN�Z4�CK=��i��c��ڒ'���e�Ŝ�i�����\<�S	���#�P-���|����9>�6���м4�m�ol!`xGK�C1�u=�B�T������&�����aG�	Z[��⫂��H����Ӵ3��=b��7�'�v�K6!.pt����zŞz�E�ʄ�v͡}����|���N��!x��n��JH���s�3M�l'O��^�&�<.^����p7���R���5#��:�f�=������������Wѭ�>�}��˯�[fl��V�� ��Xd$�8�O��rK�>�~�?$pU�������
�?66a�ϝ��M���Z����m�+W���KX�(��Q�+�G�,Ӗ��/�?�o�<NjE|��-�luE}!E?����w�:%����M�!p>$���EE�G�Y=_�F�~��L��<Qʴ�f�D��׻(�͔��)<G�
@�)�(p?�OU>�Z��	^k�Qʟ\t�	ߑ�څ��#4:"�+<e�Y�̈C�B���6�����������?���i�-o�����y�Ҏ��GOBLڍ���&Z�4��U Z��`",	3i�>�GҐ'mDh��w���aGn�Ʈ�z��� �2�4%�F����Ӥ��±��#O5�Ci�z/���r�4�W��'��3�� ��KVG�|t���� �2Zi�c9� �c�KC�Qi$TL�<�U8 ���,B+���3���SY@��x�.9���bg�v�� I]�d�=�2�=����,�,Z�l�!�4O�����1$��^�XVXt.H�S�g`��~g�&)�M~) ���#m 6�P�l�X^)+��|20x1*�lJ�`���e�O�-��^��ƣ�D�<���Ay�.)O��Q,��/��v��e{�� �}���8L�W�We$�Q�����:��F��$�z�M�K��@���Rua��`ww��.x�)��.�5q�ve�S݅�(&-��P�,��F�jܤ���H ��l(C�8��*�
y���@��h<X%Zv�8��mA���Ӟ|��mυI��BXF��y_1;e5�j'9�|���A:,�P����������5�#�Vk�_�fB-�P	<�W�&�4�"��c�U>� ̨*��
'����3�2�O���v]�JqѮ��Q� �M;��ٟ����Mda��Ȁ����Vի�%l�l�n��Z��-����vvm}s���֮�5��Q�L�9���^���wx���N���+�yzim�^Bx�=�b��v��g_�㯝�n��������n{�����)��K���i�L{��`J&xR���+���$�\��P��~V�o�Yʲ]�(@1	�((��Xc T��)o8�@�Z}���Q��4�V4"#��p�^E��ܞ�~E�5Q*��1�Ss��q�h���dJ��;��h����F4����H�vp*�q��G@t�B�h�Ur��#�@-䶠ÁL�7WP�j5�臙PWE�N52n4���;��d��l-��˒�n'g�|k(	�$p^�L�;x)^�R*�WY{�ت�֟>bO/��U�X1s?<YtQ���R�=��ia�<�{���,�\Zg`*IP��&*U���I��]ط`?��م1:(b���8�Ya�BQ"6i.8)�x�� ��~�NӮۍ��l}�����e�(���U� ��?E���B�~��Ej��
q`Z�����(>����O �4�=��.A �j��A��'�hsX�N�]���Iq)�����7��ꢽH�c��hnL��yJ�P�
�j9�B����:�.j��-F
�T��| !���e�t�˦\��0����e����w;�K�����p;/Q*%| r����5MbOIsf�Fբ��}�~��}�������}�7��-������bi�[ry��8	�·%�^�?��rdy*ʄ,Y�\q��#L�LV�:�\�d�[����]���,A[Tor�CB���P��Y�O-���v;�c��)߷֡�b�lm\d-�+�g�3�o~kx��@��B���yAM¡+W��*�^C��?<��e�~��b��p����w��CJ&mh*�[�{dqK����JU�\BIՠuQ4���#,�	�o�O��B���.�梊�E���E@�'�c\� �������4�~s����Ǯ�_�䝶�晠}��7?e���S65?o�Ř�����w��|,%,��Y�s��ڠ?����U693���+g�]o�������_�o��V�/Pߖ[�v��i'�p
���͵-�[�d�����ݿ����c9s�ʿ����<aم;�����>a��s��,	%�a�~�yrV"�}��$�'��s־p�F��S�P��/�3_!J�@F�w��C���C�x���<���ʀ"����qx�V1w�X�h���}�Z��yv�[	��<3��Q��#�� �}@��sݡ`K ɗOsт���z�O�(�*l��pm����W��Q!�+ʠ�T�y��e���S��F
^�H:��oc<	��jnnq�]w��v��;{� �;�����j�ɪ���*x���^�`��/��Ob����|�^�.��N:N)�S��ò�iH!Gé;�x�J�qj@ռ Ș��4����Ҷ���]}�!;|�����4����n+�k����AH4/�+;ߐ$� l�rYy�A��u%�$�4�)A��q:Ǘ�BL�c��Q�w���k�6jWd�ל�D�,4T%-����h�ڌT�@��y�����A��Ɋbp1K��\4j�
$-D��V��ӇtE�h�>�a%�7�3
�4īC"����C�ZԞ>�P�T7�����	���"uҐ������n�`����{'ǳ��z�^x�IK ���o�hΚς����ʧR�q�7�����4ܱ��ᾗ�\έu	%ma#�LLU$��n�a�0�=��}�K�[(�`k���R�+J��h�-��z�R�$� �.x����Eъ�\i%���I��u��H������9 �%�} �a�n����3F M44���Z�\�P�-bX������3�`n���{�E-VH-)bT
�+�Y͉����`x��8�u�W�9;�V��"0G�j#���������F@��;x�S
�!e$S� 	A 3�i��+���@;n��*����5�����5�<򻒐�r����$�4�LN�P}*�`���`����Z='�"��hb�kq���=a��Ͻ�~�Ǯ7mN�v0������˾���mv�~���H�~�K`''����B
�Cx63��~��6�x3mssv���3��ւ��It���QU��t!0J1�Hp����C������Vw����?�����>�寷AjfLh���G@�6`0x����������w�r����O�4�?%�Y�;`Y+�*!�κ+:�ҡ�d�^�1�7a�ՠߥ�II�B5�����W�:���O}�9��ҷuhY*�+��T���J��w�i�����O�)Z���Ͷ����9ڤ��-��R��O����Xu� ���@�ȗP��-���|6EK
�'�@#?QYt<Oaiw��cc�Ӏ��׾����ؙSg��+G-/�wݔ��_��^��>�k���j�i��p�ί7Ў��&�����҄ZR�����¼3�ݝ+h�:�@o>��U��6�M#��X����Eњu�V��>b冝��lgN�������ɐ�f��U�Z�h+�s,��60��VV�WoZ�T�B��R��C{#�q;�;����ƚU6֭Qڶ]λ�kV��.��J�U�-ں|�m���.�ᭊmm�1�;��]����\�d�-�b�dj�  ��IDAT�KV]_�~AIy}�����U�(���pl]X���.�\���>M��k�z�N�}4�0H�.S�a�խk�����W�^�Z�]����@���5�6)g�6/]��@v��Q�rm�U.���S|S�N����n��6�n_Z����س߱�/�d[���*֡˧NѶM�6l���v��籺NZ�z\<}��C�8J���m����֣��'m,��;��և6Ο�����k�q�,�p���K����e��� VN��X��:�Ϥ�\X�WN��]��҂5*���Z @�G0Ɋl�|���1���[���vfZṜTe�f=���X��3I+�=�u2Y�Zuת��!��\�vW�ؠ��E�E����
(5�=�m��u�=K��y��>�̺��j���<VH�v�!����g'���R��d�Jg^�ri؅���5��H�^����'��M76�������mhcqzښ�up�<��h�8`��xߦ�E+fb����U��Ҳoc�1��J�d.m�����:��Zh%�.�].MO��geh-���ة�da�>�E�tf��𰱹
���B�`��B(� ѮU���M�ʚ`-��v�`�k������w��E:�� G����W��7�?�4��x���<��/}W���1P~z�zѼmcA�mW|hNG�>�յ2��BU!�bs�el����YV@�

#����q=�mHsL(�a]SH���o�ݦ����J¥��=��(P��Ω��[
^̚��Xܲ��|� ��ąL��d�HQC��eF�~,�lqO����,,p�g�ד�'�	I����k<��R��PrWpS�J5vf���@AF�����Vu�U��Е�>P��Cs�H!���*�i�ʑ%�z�R�3)����J�zí7��xX�� ���?��lAG*R
�=)��zڡ\� !~"��%p��C�
2 {)���8[�ٵ-�U�����s��G-V�$�0 �k�4^q	R��?�*����(��{Y<v	�Uc�jN�ɟJ��V�iXK�/M!��aN���)p��Vku;�Dަ�y���y����w�i?������'������}������}����~�C\��cgs>��x��U+�����d+��D��E{��Q��������%D��G�L���LA��\���8�0\md9�@.&�X�!����%�S��>�+[�]BCmX!�C{F�)�A���`;�q�*��:�Ss&�	k5#Ks�c�"�mK��;R�� f9(�L1b��L&[[�b�cy�T��C\�����A��&y �9B�MK���c᷊@D9�V^������sGm}�8�����������tA��E�"S�/��&�b�-4�v�$���U���KO٣�gNEH����S�~�5[G0��=@h�66�{um��i��9� ǐ-��,�V���-�L�88�G�D�u���9�BZ{��v`z���wv,Fha{�~�O�L>e��pݭZ����A�����_��g�dXb��,�چ٣����`�[���T�Gy��<O��:<?a��iwjW?vwVmP#�C9�ύ���L¬Y���C?5�i�2O;f�)�<��(,�� ��XU)�va,K[�o<���e|�ó�CN�6�s4-�҆n���:�k��j�ffm��4�hӭ]p���_�2�O�g�r<��~᭎\��920�%�\�C�3�S{{��(*�H��h���M�k$e��o�|��7`��=����\�� ��viC�+kC�WI��99��+�SW��c�#�©Y�'��-Z��@�ŭ��[/2�u7��7i�����Ʀgo����+h��%K��"+ �&,�� �)���u"ykGu.z��xz�V��J�j5?&|ȱ^C���%d"��S�a8O��%�F�ϸ�r�A�U�VBJ)�D0h����D#�lX����M	تf�\��9>"7�vA%aHx��5j����Zk���r��q�$u��|94g�C�J��=�`O�`��PF�u8�\��ҋ�?�j�������*n��-���/����¼]	�沶�oѧQz(�-~@�Bc$o�� =��E��"ű��n��h�[I��߈0t!O�o���$�<�$�I��c7�1)�DZc����w_n�L��Z�X]��%KT��wM�o�f��Kb��&
����|-�4����}�G��I�Q�)WZ��܌M�ͺK�T��94qm��=��0�'��)C�A�a>"�L����{}�U�m����#m���(�FB�;�*$���N:�х�icŨ��)|Tp��0~'3X�.�;�M16��eB�E�,f�6V�R���Z��9�6L}�-L#�pK�І�3�&�����֨-�+0M�ɏ�29�0�h�_��Yْ�6��&`,����w��M��Q@^�_�U����X�Ў����i5��8L3C�9�q��)ԑ�`	�M��e;z�Y{��G�c�'ZLr����k���Od׆�]��i���l����l̊�<�
H��F)� Nu�-?��\&!�<,%'�@Ղ_��'�9�D��|dO�ְ��H[�+ֶ��8̰�����~�zi�o�m63]D�L'mr�!���!`���E-�����B,B�4�Ӓ�
Q/�N��i��K��9���X��|Ʒ7�ˇ���Hت�4J��g�s��2�vm��A]�>V,Ƭ ^*��ڐF)P��(ml67`����N�0#hB��b�/#7����X��Q��@/B�]$��y�#W$�X�fn� �Bት�oǦ���t
�Ćb��Y.+<�ف}c6��K	OQ8"�/����A]�6X��mom�K���(e<4���u����G�9� �������%8�	�¬��z0�ְiX�o͟k�W�Rrɢ��4��<*��x먴Vq�6@�Cq�%)W���KڅKu�Cv�S����`�~4������1�|��_W�ut���4�fOv�@Y�o^����@wd	x
�*��%�t-[S������(J�xuS����������Ќ��%��hNU{��>ť�+���n�	䈌5�B��SX~'JZr�yUyz�h*4DsE��)ɩ��Z��l��ъ��4�B澄�����Lm�V�h����̤����%h��ʔ{���V��+/�׎���<�=����ķ�o|�~��+��}_����ůp|վ��/�sO=ig_?n�4�|�VΜ����S�>o�X[�g�V�hM,��K�lk�4����Ӷ���-�+X?%����v��Q[;s�6Ο���^�ܵ��΅�V^9k���~���$�:͒5kV�����{;��Z�@~�m�S@��'b%4<*�a��%4�u�<�B���F�"����|FP�*[��Z��xSՂ����cY�5̄�_ټd��e�V�,�&}P�Y���UU�ms"�[�X�|�<o`A�a����Cؚ�Ԣ#-��ܡ�h.W�����6�,��ל]&��y���h��{��g,�7���fe�g�&]��a��e5��mC*}��V8�eIB��q�0i)v_�G�ZԂ�0�3��j%��$4�Ҫ���!V���War��<�Y��A׆�Z5�~`08i�K��.ֵ�P��V�K`"�C=��7�7h>ASw� �Hc�����]f \�u�ͺF`w!�.Q�M"�\�\(|mֲ�A��f{)�T�PP��^�/��5�[QdP���U���cע�!���چ�Ш�����G�%L;ȧA@K�K��N��Ft����	i4����V�h1J���fѤ��� �u(fH^!,7�ڏB@�4/-W�$|G�֚�ˉ�ɩ?��S\+�p�F�������o��Щ�zP�5��n�`��1����9h���/;�+�\ަ���;��lw�K�-i���*�:�(/?�C�;q����4�Y.Ehw,��"0a��v+0��6u��Ĭ����P�&@�9<��W��HA��9������<o<�����>�	)z�O��	��ֺ����t}D*�r�'Zĥ��M�bIsv��bn;��Ń$��ă�P?_��z~���V����ӟ�D�J�n�<��-ovm|r��֨;��d�t�"^u�ƙ~�l��,�����.�Jg}Y����n��� 7f��*�����-j̷�֝���v�&q��}끇���i'N�x�N�Ν<eg����3v�W��i�����?e��UJk�~��n��෸�emV�� Ah�v7�]Q1�{$bm�$�vy����E��C-���U+o.���Է,���J�s���S�o:�
y"L�X"�L�F}��+�Q�A�V7^h���`�����>H���s�̣��h{�mۡ>-�6�vۅS��vQP:������.�k��@��S�G�f� � �i_����b��������F	�!PT�%�Dz�ĵO�T�Vޥ��������0wZvȂj��+��X<�$u.A�(A��K����'m	�jۗ�{Ҟx��5,�)���f��G�+��h��V�f�y��]�]��Tf�������3�\6���x!��E���y�8mU��f�����3���B�ՉZ�0c5�Ҳ�t&i�.\Ě���`�Qn��<yU�5_\E��G����NB~�t�ri�6� k-!7�A�=�hC�Μv��"�&��Rc�C�[F���6v���$T��X1�u(�v��
�_C_�%tN񽘬�{2۸���'�I� @� Hg��Z^��±�]�6�����Ɗvqu�PF(i){�~�����6���T�Ϝg�.h"�R�"6��ė/��*���^E&��|�`��^w׮=8f��*��EJ�677�s������1����@˹b�v�fg�=����sh����I_��U�:$�vQD�(�MQ���y�
��2�.O!���;5��l6�oh�o�����u��v�=wю.x�.�������Kg@�i�J�|�쌔�u^��`��4?��(M�}r�5���N"�7\�M~�Iw��*������I���t���M���$�Q";x�Y?0A��#tzA.H�/���"�u��.^ ~R�DS_��'���Ց=�Óe�[䞤1?���ϫ���8��4�I�J�S����ܒ�j��3���,�*~��>�iY`w�(g�Ե��"R3��P�:Rc�0a*/�*-J���f�V*���K�E*k
�jjq Q���-ʳV^�����@Ph����F�����rì�O�%���㖃 �h�㙄M0y���}36�FA�B:d�ŔM���c)�)wqv�b!��,G3�Dm,���<ϧ}��,�g4�FlM_�<7���������M��5�WǜV����jNb�@IK)��АLJ�к5�2?[�a�6��<f<mŊ�%{tx�#�hhj�&�h3Z��@����Mй	�����;%��+�0)5rީ#t�w�Jz�X&���<�1Ťi!x�����@
	�)B��!�<Z?H�a��'�S��h�-<耀a���B���B*�P~�ڜQ�|#�z|>9ՊQiY�����'8��V`�R�.�V����G��w�-�������<V��tA؁��T�	BC�f�zW+(#]�&��8�LV[��0��RC�($�����HvM=�����!ߤXBX�v�&�0�N,E�| �ȒłD�ɏ�/�5�����8b������
�s���f�qg�U$�"h���8̯M�r�\=ZX'(=z���_���9�S~��Qf(�p���<뻃�4j-w6V�ta��g��<�uha�T1M��0��e�c�\]74/%A�ḒE�)`NPw�6


�nY�N���u�����a@�Z+�+�!�6����NV��h7���C�k��{�����;�|CC����9{ۭ�(��R�j�lzvή��z��~�>��{�����?7c7�p�n�z�n�~���-G����~���w�u��7	}���Ó����f���箫�}��>��w�?2�Q����z���ٻ�y����:���C��0f�O�M7�;n�֮�
~]h�B����e�<�
m��ߣ�U�q�7��T�$b�#��CzHW�-�׎���� ���B���]�=J����{���g���-�Fbl����"�'.yi�NR�q)��lZ,�(�be�"|BJJJVH�@���$�&���J���6�V�8��Rתz�r�kM��\��H�Ӵ9p�g�-��\�I�{޲h�A�B��֠E=w�b����eO�ִ����h�{A�FFm�L���ZN-��B��AP!x�����$*b�!
1lIa�ѻ��
�����a)+��X�~�������i,t3UK��n��9_���%���X@*N߳Ͻ�{*ɼ�_Xpƛ��Me�0���c��D$i��͢Ah�H�LZ]Y'�X5���C����LƁ`?u�mmm#�����633�Wt�珝&qK'��)g^�	�w���ًy��+�8Z����s��S����N-2�Cc�|��'�h70�A�'�7��ڬj�Պ<pM6듹�k��B��e���S�SV(�(_:��hR0��=3{��ǭ^��B۲���yTH�+`�a�L���_�N�v�W:M�Lч=;����^�.�y��-����i,���ML�ҡ�Lq_��m�ZN�W��\��T��;w��eb+&�����n�(%[h?�����}�;+�J^��BoAk�KY�UC�Ӱ#`I���lVC*և���Uh؊�_�,m�kV?��n�~�*<�NS��R���)��긤�j<Uȶ����('�N��v"`�Q#H��rw�vU���
��$ZF�0L/����"�4+%��} �d&m��X�~�{(:Z���;Mw�1h�r�)'ն
�za�r ��V�M$Ђ���Qh�NBqk�p��]<Bߥ�8����w|Z��$���;7:�YV�|�4_�}�s�Si�\Je�/��݋���Ig��.�\�7�<;p0)
r���֨�Y����߸�~�n f�=�W��J����O`%��#�4T�$Gy���h�O�DCÚ\�H����-X��V��
He$7$�W�ZP�,�2����N���)���|�9������"R@ȸ�e�8��V�	:�v��SN�Z4��8��ɇp$!�'|s��a�aB} �z$+�[�_}S���\�Õ$+T���=�	d�����\\޻ԟ�d������t6��	χ�44�}X�Yـ��e���Bư��91���u#}�*�w�G��°�(���,�,Q�l��P�SX����o��ν���./�{����~�mVhc1���������o�W�bz�՗��>\�!����@%<$��\�k��|�$���5~݅�j|UXS���6��f0Y-���6���tV����ۏ|���� A�ZUy����o �B�?�xeqJ �B�IK�ݝ��*�d�*~�&<�h�I��c�j�榘==���M1#,@,Du�v-V�U�_$����5G�qgEK���FeU���V����E� a�N���1,j5!<L6�9�����0Oi�;�)
#�K���k֥
�4oEXО*L����')��|�b���dM(T�"5�g������K@k8R{�i#�LD��Lg|X�L}�-)EL���7k�̹<�J���O� ���U��ǰī�@��`��klk�N���G����J�H� �F��qVH��]�<(>f����~���>����o�#CsA �� u�+Pv�v���}�2��N��%�1����ݒ�}�e3*��3,A��v<��R��n-T��2ð`�A)�FAM��j�|Ġ[_]K�)l���O��a}�}F�������!�����bi)����<[MᏴsu�ea�dš�橰y��������J�G�"Q�h�P�Чک]�e5��"�h��� ��};E��0�u�����gk
� ,�|j9�'�p��1�j[)9�s��H�0��!�s((��_�G�D���V�bT lAA�Ri�V�j8?�8e��������e�:i����]x�$xsXr!�����`#d�0�"���o(ba)��_�D���x�00}�x��C���7�
�P��iZG�L���?c��w�f�ɛ�b7�k�j�����o���-I�7�ڃ��KRDeh��I��L�T֞�f��7�I^y�W/�����{r�Iੲ{�������&��a�4jk�W6m,�@���55��M���T)'�6 >�4���Or��L/m�
`�@N�O#�n��Ξ8ik��o�w���o|�Z>���=��[�B3��G
'�"V�,Mj�~�C��d�h��������Χ`��i	o���P��ȓGi}ŻW���Ʉ�qv�����m�ܫ�~���jK ���ַ^�ncc)(�5h�,rM�ԩ�0���.�����k�ZHQ.��[S`V�h�cm�!39�;9�(���L�}C��Ea	����$"��ӥ�ԵZT��!ЄG�P�ғ��R�2e�jsbS`ia�ғt��Z3�H�_���s�&\����Rk�9�������V��C+U�4�Cwy�����5�м߀24���"���js}�!j@��
9�U��n	͵�BRm�!ȴ���&B��NE���NB5�;YM�XH0$:R#b�;%�؞�( ���}Ʊ�����pl۞{��������ձ	��:o`q����^�2WV����7֛UJ� �Bm\�я�V�:g��e�
V�����6ʎ�ho���j��K>�+Vٹ`1��b%fLJH�ƋL����+��#T��s�5���!�m��k�\B9Ci���:0h��y,�"�X�h����[k��݆���&��άY�Y����{�_e_���	W�;��]��<��Y���Z���v`�(0��3vW�E-�����6���)_���	۾��σˡ_�v�uD�61�^Y>ԳZ�0NkAL�iW�R8�臲PTL���U�s�v�S�h�s/a!W�c��v����6 �"�˫���L������5ā����k���~��`	=k�,�P����#�$Y�Е4��X��d�R]Y�ƒ�c��4!��:%!$EQ��ʒ%&�V+���K��>��?|�^=����"B���^e��K�(��=m����U��F����u�w���J�`��@�V�P�������%|��
\�P]�ߺp���j����Kٻ��OI��~�m��;:�g�oNz�ʥ��T��=���O<KRQ#|n%�,��-�!E@�����#�F
N�$V�r���&����.m��\:(4,�ٹY��,�<^�Ӱ�«[-ѩZ�7��>�Ք��{���va����|�emu�W�h/*��{߅|*�3s����#)�cS$I`�I�je�%؛k�B�+�H%�$ ��lin�J�ˠNM2j.m�cO����~���J����Mq3똿ۻ-{��Y�����4?��N	��5�x���{���<����i8R��>uz�Ο_E �m�TG�K�U�)V۶*M�ݎmb靻�a�/n������P;�f��]u�;çak7�v�҆k���W4e��l�k'��.S��E��ϣ(����׎_��;j+|����r���is��$�[՞}�%;}�,�׵<Lsfj�>H�W�v�:����Ͽl�;u��c�k��Q�T��S��K'����E[Z���Q?4q����u{��(���7÷�kdscׇ8e���N�"�`� L����=��s��K����>_P��$]�����X�O�x���'c�IpC�8S���{�����Q�Ȧ�
3vx���,V�+(�&k69.%*>e��1�ø�/��4O��R�X���ٴ뮞���6�����Z;�v��MLxL�N}�n�f�~�C7�G�s�}���;����#�f`�-;���>U
[OrK�Y��I��WA���O�m������-W��ل-Χ�#3vp)oW�/�-�� ����KOZ&�C���<��CAR��-ΌYm{�:��b-Z{�n�v�n�v�n�~��Me��qѪ�k��2R�������ԍ�&��{���G��{�}��o�w�u����#�0]��l����>w�:��|Z[v���~Â}��w؏|�v���a���;�����q��;�P��Ɉ]���O�t>b[˯[��0����(V���U�Gm�s�n��l*E�nQ���rÄ-����X�ξ~<��"

34;3��V�E[%[��wA��K'��딅U���F	
m7���-� ��x;C��Ɯ�9�[�X��T,IE��n�.��c���o?k�5���ժU�-�����o(�򡼶�rz�.���~������
�0b�
��c�W�/)Tx�6��4|N�p��29Y��6ʌ���E��BrkM�Y�]\(8�>{�
�J�ߜ��~O�v�����;���7:��{���\��9p3��J��F�~(/��/�g�F�BF���(�o�R����%v����P�V)k���dɥ�njZ(�auE�Q��z}�ws辠K��jQQkx�\53;k�۾zW���s.�R(�Ѡ�AFf� (�R ��涪��$�4��f9�X�U
�)i�@���.%�x������#j�_��Ni��{�
�z�i{��o��glb���v�A��0����v_h���㶼�b[[;#啗��l��ާ��.��9;��+���Y���n����ڶa�=v�U�q�������OL�۾�f�Jhӯ�;k�Bб��-��#�Ds(@p
ػk��0�){���'��������A(���a{����^��������c����vo��|���'�v+�曏�x>e�L�֛a�����G�_��5 ��n�����w�敹,��������_�ٳg����>d���w���=��}��_^NMه>�^�V�e}/��R������|����F��v���]�y�������o=��-:h�ȇ���>��r�R�*X��������r�n�Bvם����u�jN�8i�{ݞ|��¬>���Ȓ�gb��3O����ӗZVjk���Ua3�x����r͞����[�|7������|��v>�E'�b\QV�I�vV��������Ų����>�)�Fʦ1�隽�}�c��{ڒ*�ŉ�X��.�c�룯��/~a�VN,[��M2�V�La5`�������;�k��]����ZB���Y�_�b�6�=b�.���ug���m�]�o�*�GmmAq��q��������N��y�]:�"6�.��by����e;u���h��;l,�� ��b�X�r�^;��l�gJ'm����S�����&�ᖃvˍ��t=�V�*�:�m��k<�n�o���h��o���)���o���8�P�W���~�.�#��"�i~,��ضw�q�~��m��q�۴��5���Z}��B��/LYs!�������>�(�U���]w������k�_������o|�	��PrQ�5o/evqa�G�z�U{��b���E��XrM�zX���N�\��R���n+<���/-l{�=��w�W�>����#��C?j�X�^�ڣ�=�����~
�]�9mJ{���l�b׶�}�L8�ѕ1��f3i�E��Y[=��&�0p`.�L���I?$:�W�%�a��s?;NIL��M��p�ɝ�IW�F�5��.�� �t�^�_ߝ��>H������(0=x ��G�����#�K���m�"����!����e�6����/�-���$�F¦��4��XNX�� C	Z��M�+�Z��D~�W?�i��U�a��C/�j%b��Y$a���WAv2E[�T8�za��B+#�OSc�%m�Ѓ����J��U%�!�z+
$h�hNrJN�$��N�Mҭ�H!?!,��e���k�b�� n[Xu�?�}�sߴG�:n�b5�&�V#dɱkGs��w��g�p�=񝣶�&61w���Eg�'myu��I;��Y���Ԣ姗ly�l��V���;0姞=j�v�cY���m�����)y;fŞ{F�+�z�b�zض�!��eӶ[��+�����v���i�\��'mz������#�?kOk_���Y��]����h����c�`�n_��{��Svq�QE��Xq�������y�}�'���?j�Ϯ�Ns?;ec�QBH�kٟ��߰O^��S��.2K6�m���g����W��')�-Z;���u��C����g���/������3�~��ɗ���=����>��W��i;~f�Xn���i{⹓���s�{�%�}�^� ��m���������=��Q{�U��p9�Y\��7c���q� j1�_�?go�)gz����_{ �1��1�3'��[�Q����ڵKYK�dΣU?��6
]�r��;o��~����tȦ2b3�j�	C��X����^(���^���~��NO��Ug�g�}��w��V�R?�F�U�X�)2�E�#Z�V��w�#��_\��}�ʡ}V[X���*�څ�����k���˟�[���`�9��A}`O��r��(����V�?�?m�`�N������V��7!+��RvÑ9���sN���[o��~��9��`���E�UEIBEvX���< n`�`A�#�[ZC�<k�ǿ�g��{o�;�L�-���O��^Y����TΊ���F�J�O|���fO�k�($[%{��IKB3[�mޝ���);��7�l�8w�6�xQ�N�������c��?��=��);qf�j�V�{셳V��ҥ������i;�R��F�*�){��V������u�º�G
3��oO�\�2��,^m�>���O����a/�X��M+�66s��;��',36��q��|��Ҿ8�`}LN�p��1�6䦒)θb����NO���3֕�Rމ5��Wj5�VFy�p����3������G?֔�B�4|���� e9*���XT^�/���Ny�]	�ī5_ga0H�����꾄����{���� �|��ګ����i�Y;m�1�O��.���Q;r�]�t�v�� �0�؁��o����M7����Z\�x��-�E	Jh?<J;������c�k�:�[?�?U�d�c�h
��Y�h�k�'�(��6���N T�P�H�{D����� �㤱��ci��r�»Z4��175�%mA�C���&��#��e[������|�2�T+�4i��[��r!�� m���J;i�;}����A蔻i[����X��I,�Lt���%,�;��M���	�V,=�F3n�h�]��,өB�K� ���]�����歗��V�H�yk�Ƭ���j�6QZ��5Y�!�s+5��G �n7��f',q�cw�k�n�"�q;��ˁ��p�e���u�C9M'�U���&�Y�:M� ;oU,��~�ꡂ���鵖�T�܃��;=��m���F̎#�_>�e�<�>��q���K�fx'b'.V��jݖ��V�?��6�_ӮOo��Ͼn�8�/��Bi��m�g�ϤEx=��9{��%{}�eg7;0�ԅp���D�ٵK0���a&�0�K���_2�^���9�&fQ��u���}c���i����8��0�����z���y�d1�jܯ5{n�Ukm�3;�d��y�a@���$�d�2���k���?h��Cg�`ph�9��;�=5�#��˿�7�;n���
L�j?�Cﳏ~�f�D3%��IZ"*�O3�Z���'���v���������.����[�!U��Ӳ]8s���}w�������l��R��e�jK�D�D(�]0�c?�^���V���=���G1����je�����]��~�g~��0�:��D {زHg||��(-�h��jZ�"w���Q|{�:�������/���e�p����KE�j�m�Uó����	+*���D�⩄U-6lQn�~�d�Zri��Z�/A�����&���^��[I�s̶:id�}ud>��/Y��lg��������Zl�*!�`	)����6�)%�܋��Mڲ孛_�^~��|�r�zY����Ak��W�F���q��F�jX�Z�b(m���r��o��4�I?x�ig9�k~NC����B�a
\��4��$f\�H����HY�� ��C��vuHj��`�^��{�!�L�
&5JQ��L�y'XF2*s�(� ���x���TZ�E��m�("��C�qUg�����?���5+ժϟj��"l�-u跊a�����C� ��M�/�A� ����'L~�o�,�?�ԧ��-+�c�Q�ZM���v�Ee���SR��~��h����jh*���L�@��!��Bٓp����R?@ڼ"N�F���'HZ1�h.�"o`5-\ ��E��yLт�6����ؔ��k��.��[�֤�  ��p���8����9-G�*�Q�|#D��,�:H��C�V?j,9��[�2:�����)�7[�z-$��X�� l���B	�Z�9
�D)�_/K+�ȣ���O�7yD�>����d� �Je5U�2@\�H�@X�d�\D���t^�c&�/�ҥ[p�@��'�=�8kۣ߻�p�a�1<�&-%M�IVfGN���{��mf�?Xhub�۬՘��F��\�`]gC���CBB����;/B�zq_ɩ%ɵʎŀkJ}�����Ӧ�3�<�5��=��-�Q$Oh�!�X����W�lA{���W�����MMM�/��q���V��_ްǿs�^zu�^>�aO<��EC�ݿ.PN:�	<k���ɓ����!�������A��n�N.���V�^9�m�|�E;}iǲŢŒ���};��}��S�[�P�)�ɤ���©��ȡ��̏��ͣhR�>Sz�;��ǟ�6J"%K��و��������7ц`�a[^o؅��?�e+�M�����r��o��Nѷ��}_G�O�;�~�[q�ñ�]\^�u�s���������K���S��R��w��n�}�?c�O��m��b���0mۭ�}�O�K�����>� �J�ĸ������y���F�����_�W�l� �ꃟ�ށml�;O�җ=�Cj̪��;���b�m�.I�P�w��0�ѧ��e�s?BZ~�=p
³�ml):�V�B��v�
�{��{6�wL��Y|�[����;A[���VƳ�G�@{ʯr�T�!8��ÃN���*�߷��U_0�1h_|@{^ H���DJpE�j�'Y�	�g�^(��d��SC�A,K�̔��{�f�����Ą�>�|��7����G���C?����	�RҲ�c��Ӛ�d�B��h�I%P>��'_���h�^#5Zl��%�D�K��㠝�NYZ���~m�X� 4}_k͆�a�MLNb�U�LǺm�7��w(xt�i*�v�����Z�
S�@P�m�ݏ��VO��x&Grj¥��GF	�)��ъ�kY�o�U�M���ϸ&_@4^ڊ&5�YN�rhm��MY�L �h[{��6�ڱY���$�%�Il�|���b����qa,_#!,�KPQ1 ��)���!�Ah����W����!�tZ浐9�yHSU u�"��Ѽ\��u@�k;BǨsR���vh�O�Cg�jS��s���EL��!&�r_��nJ��X;k
�'��C< @2��h].�`}[�+�@�[�o�)���6rLTi����7h�7
�I������=�E]*74ڢ��ZN���c�:&3����M"���P��S�a�\[��*�~��j�`��Xb�)��w��f����=��Q[oP��]�����m���΂(cO?�=��w��{�a��M��)<���|��?�����^�ǟ;i_}�	�a�s�X1.��M��c/xt����?iE ����W��m���������~���C��w���H�`sXAi�Sh��*����O�EB;Vοjָh������Ö��e�Q�x�5�?~������v��p(� ���?�6;����=�����o��߶���c���Nأ�=}j��e�1t�43��G_�#W����.wc�@���t�~�w�о�oؗ����W�i_����G���}��^������/ث�����뮲��p+x�ڳ�}�);��kũ��\��99��1���o��Xp_߬������h[��U/-��T�QvA~�C>F=[-*iv:�-���F���d%M�;�
���� ����)���w�v���7S�x�8J��򨀓
�(촥�F(t�XA��)a��4���(eQu�i�V�qf��R���(�M��V����|.�5�� @����%R�\G���������k����Qx�"��ͮV�B_����;N�4���~�
I�%樲U������Cp_�Y[�H�j�~��-c ���OR�E�y�a "@ݿ�ʥJ��Ji����]|R���"�UѾ��g��;�P�hm�Z��|͈`�D7�̴mŶ8>��+�b�w�M�\�)оڦ���&	'�=�<n��V�(c�h�EvU��z+@k�SH�U��ǨC=�%�4=m�z�ӜK��p^Mvҡ����,*�҆ �>D+`�yS�����a�z.�W���(�p�ϥN�X���0V�H�G �v��6��Ga�^�Δ��M"t��\�H�)i٬��зnM�)Q�m���|a��:�MGˊVDu���zt.��D�Qt	^	
�U;�
M�"�kO=�͹#?0ֆ��W��V1�	]���d��w�
  $�p�&�)��B�ȱWLR{��yȢ���oMB^*������pC�-�	����[�x'�ݙ�5W$<�U�C��׮澗*�h�X�S-�A9��+�E9���!�xAE�=_�,B���0T�I�2�㪃�a�0�ږ5iWbmү�?���t�4}6fŹ�/����vf#f��_�?��Q{������=�����
3��T��FF���'�cgl�ԳJ7g��[l���?����{�y��r�|z�>��'��a��V��. x��7~����r����Za��_����?�cgKֆ)W�[/�ʑ���Nž��Q;���i۟}�y����"�<e�7�0����v��9{��W��K�Vw���H�7����k�}��}�0n퓟�������������j���{띷�I+����rv��7؁}��EC�b�f�g}5�+tY)sI0D�_[�XF_`�
�p��:�Cn�I�Ҩ�"�hᑂ4+PC$�]�}�D�����:�2)Ƙ�����-L8�I1�(��1H��0����Xc�"8����NZ���B�XWM�Y��-Ǔ�^q(�Z�L'M;Ӄ�V��Nc��\9KS(���^�;�Y*�]NAq�B���ɪ���:U�Yal�E�	� �����8X�����N��K�Y�����L<Iϡ�0�ƅ,;���,�!k���2);r�5@m�Պ(<�y5�zR�/U���ѢEEO�4��ݪ'�-�B���N�d� �<��RՇ43�6���_���mahiHS~{���EL�΋�r����a��
�U~�do����e�����?�����v�>�ֱ�z�.�`�T�լ��N��X
�zA�NS֘\
�Ѓ��O���1M���S��ڿ���
�끈����h��T�D�Vh"~l,��ݵK��`�
K�Ɠ�M@T0��,o���աʒ���5�I��*{��ר[��5��
�PMꓣ>ڵ��+_&�1�-KK%SX�uJT�;�^Q�rV�w�E�.���������w_P������� �H*W��Tx1L�ݕ�V���!x��06	!H4;3kk�O��S��NML�r�m�*�ze���(R�U���FV,<�۩�.,����K$��s��|�#��H	��s����;V��ΒWk�Y�W�j,>�Pѻ���V�نICP��4V��E������J�c�Ѯ�ͺ6)�?��]�RG�]ɥ@C;�iT�ߌ�L��oU��K�,��62=�ʛ}�Co�ix���N�ky߷�ӊc)W�2��LYŐ]�4mGs��i�+�������:��&�GQCẴ^�/|�Q�i��d�m��ED<9[[��ꥒ}��_�g�z�W��e�w��!�"0�����"VFʶ�	¬#K{�<����G��ǟ����7��iD"	j�u��@����[vǵ��oX�����?���׿x�6���[:h�x:�:p�	A�_�/��K��SO����>����������6=�w�u��x�A�"M%�pr[�{67�w����w�-�����^����;��CKv��ۿ4k��v=̤f�_?�Y�������f��5.�t\���Ţ�B	�6ک ���]�/m7_3>��@�_~�1�������liQzS���4���(pR��6@�	�+�n�W���Ԃf��DDĤ��o>�� �h:��i J)�
^F�P|sh D�N��j&s��Ut��,)�М�2e����'�V�ܲ|m ߪV�|�͘�yO|E#@�M�_� &��F���$���Ks�>��# "А����������kQL��0�����%(�G�K�A�4؇2Qn��Z	�F	��U��G���@�!��g������"�ve�.��x��y��Ԑ��t�wNA(;����Ѣ	g�2�:�.����HB��H���;�n��݂��,C`(�-a�n�
m*.�����+DM��;H�_���G�*���r����5�������4$%�uHzJ����s�V�%�ssst,�I��uOK��C�i�HY$�V�	��
MO��������$ �ɘi[i�r\.�3�H<-�U�":i,�t��lia�
E��6@1� C�o���̀sڠ@�!N�3��[�#Ң�";07iq�"m(������9�u[��N����0��3�&
)�*P&y&ywi~��R�`��h e~�`Y��c�yi5��� CN�XD���KKsO�[H�!�����<4�3�I�D�9"j�eA�WZ�������B]�>:9-a���Y�����PN�	�(pGPf
Y;0?�d�7=E�Ϥ��ь�e����i+�4�pVN�	pamTyj�8k�6��s�J������`� �K_Dڪ�������,���߀s=,q`#��b�A��T�f�h7�oK��c;`qݍl`(0��W�J�Z�-�U�Fc�� ��Ԏ��(E�I,�y��SyhG�Y�j��A'���m�� ��#�����L!s��h�{)���
�M�`&ű��ON l����AM��R�CK��¾�l~��<PT�E]N��\�~���I����%�ҳ���MY��-.�wK�Y݂����|���y�f毷�}�XR�1���g�	����v�;nq_B8�d�/-$ӱ�Q�9���KmӲ�0is3Y��=Ł��Bt���O�Ƚ���;?a����ޚX��fqp<��bP '|���Mg��_)E���<�w�: �Bs���I�E�x=�u�A�$���*�]���
�՗�v;X�p 0a�h�G���Xes��_�QG�b��}�T��{.���H$b6M����W7W=�@ZO�ߢ�9�8Fck�V�ڰm��OP�q�A��Y޶����О�],_�|6��N.F����=��i!O�$�%L:��)��"���-�#N]�Ͳo�ۣ���+�&����G8Fa�m8�x�od16�=<3�U���T6�g�z ��������V�ʩ~8p	�}o�0��/��p�h�.�[Wm'Up����5��u����7��*��nV��P �"!^���Ϟ�GK�5*z�
N��W� E�%�#���4קm�<:*eXk���IR�)�����%e^�b���a5	,EZ��	jQ�Qd^�$�8b19�l||ܵ =�qv�}k!���-.."��)��걸S���rc�cahgt	Z��Hʉ8R'��ٹq��@U��%	gAVmF*�cr��k_0u��SK� !1x`�S�0:��$�#����:�I�ퟙ�*D
&!���v�Qj7c	;��P6D�����U�~�� �����E�nFZ���s ���>H] �9����a�8rX�E�>k��"y̍cu��i��$�!a�A�Hs�am/!p"X�bB)�Fϊ�C��S��K( ��^;�@�b:��|�IBSuP�4���/c�Ӗ���DQ)��%�{X��}��a90���I��iw�pLs��o�2I1�������,�"YLT
�V��s�4��qS�AS���4q� (�Ф�r��4�[~�Κ�>+
�$��>)����`ܕc}�St�	���u�1���q�uK�kü������x�����Q�dY�N1��H����A������/������~��7۸�EѯZZ�m�7|Ԏ?k��4mv����u&Xý�+�J��}>pzn	a>a����K���#���?����n��j��L�[4�6^>z�������@�x1�U��N��u(�ֵ��&���}�]�T�����[����#hA�m�f�lq�U)�R��I�$L�K���$���=�� ]�Î���.z|v���q}���'9��V��:JP����yoEt�]¯/W(�Q��,�/&��D��,��?(�M}��j@3@�B�D�,Z�<��oa���3qE�i�]�GQ+$�UE�4%H�x�V�ю'K�h���G�!z��>b���{��Q;�wa�Zx���I���E��]_�0pKKC{�1K��,5�K�%�7	E�)�ީ"�B1mP���I[q��F�^�L(zR��~D���>���@�hWQ�h�hP��5�����lj,��6�nk)'i��|N�;s(�:�~�Ί"��81A_P�.у.��K�~(����MMZܓB4 �nD@_Rv%��cE�œ����A�y�������˻ᵒ�,G|��*Ы��Ƥ�":}�Hc�2��]M�*���4W')l%�O�2�LWLs9���F�"b������˻!��=Z�G�����*LC^Պ��h8U %=���B������K�c���u��(Fyh赊E��]���5^�:je� ��S4ߤ�/=��*�hٰ��
 �hŐ@�ˉ��!\5n�pI�+�1q�y�F���Q�5@r����ӝ}�P-4�. uPoh�)J�`�JE�%�#k�1�`�I�Ǉ]a�4��w�C3��n�¡���<+�xP_T\�-A�J(2��
(�9h��.m���J�R�Xy�z�O2IQ�0����"�^����zrh����UN���j�꫹^Y/
l��W�4�N_hQ���^?z�.�^���1 �dݏ#s�6�V4	�,D�0=fG.!DQ�h�V�i\C�*KZ� |[_-������N��P��*Uh�5Y�꒕p���m��Lg�7�S^KXB�W�Y�U	�3I,��mD�h�M��\�>r�-6��v�������ڿ����N�9�ϵ�'V@�����h��A!�B�6�/Z��Ka��
���ٗ���o�����+20E��<�o}Ǟy�($�	��0�ڤ��*�q�|ݾ����[�z�V.mÐ4oV����Y��Kާ	�0{��<�Gy��O�e��B � C��<跬�QR� 5|�i�qm�*��h�$WJ�`%����$e�G��@�q�#�uܛ�f�9w��
���Eƀ�6}N �&�(}�q�N_��m����
=��ji�E��2䑦O'�V��q���Ku-�Q���*$)#��ط��
g�v�C5�Nj$ ����i9�G��1s�:2WsT�ȡ}�!+NA?ߘ��R�%�(Gʾ���ӊṱﵭ �f�7�E�1���%�C�w��n��ѡ�Ȥv����%����|%^�]����\]튢\ȰP]}���7
�OߥQ7� �fg����T0�B|r������C�)J�F ���� ZV����~�]ƐB¥Q��P��C�����!xS	z&:���7`��R�ow���i�/��\���9��XeT�����ӂȇLss������-��ʊi�P_Pva��ǣT[]]���ȹU˄姳����]�c�e�l[��k�GĶ�U_���.����5�Ge�K�Q�]1�d�.¸.�hY3��������7u��勾�YKb����.LJ��k�?}�m�|�R,ıUڵ��]�U�z�.^�m�l��C���nM����66��܅���ZF�������;{ጝ�x�� �\�������Vj����R�<G��4WQ��uAܥc.����ƪ�h��(��йI+�kvf���]�}���[u+sPF�Z+m�6e�!�b�:nj�A�mͥ�+�����v�����[��Z�2�[�}߷A�]X	�^�.����ȿE�u��.�@��;)C��V�f�Vw�hG|�^d&��$��e�$��3gf�OEI��9���*�n����ZTq��	;u���,o���`(�K�_�6����1��k�^ۼ4a-5m���Ғ��iJH�R��N�\�AT5��X���W��[�r���d!���0�}�Q�.�*ZXo�l����Pȿ�[!�Ů�� �VH+@��ԁ��Z�P������O|��}�%0���1�Y���b���������G_�'��5�#�=Q6基T�?���������_~�i��?��}���R��G'vi�"�ڴ��=�d84��h�c�ze��R\N�G�MN��)� =�S#7���ҧ��R5-e���p�mI�vV_jq���� �L����J���\W����a�І��Ӑ�b�j�0�=#N�I�(Ra�'�V�Sʰإ뵤XS?)mZ�!�JC�M�H����@S�_�L=��]�i�
-�!+.�������K�Q
oO!��${�C�O=�LiJCC��O��C�=�>8�]1�Y�)�U��K���^nLa���K�h][�E`E��v�!���&+N�������԰.wk�E���p�5��2�Z�������K�M�>��/�F4�آ��[��i�<�C�I�#�{*�]}�����4�o�
��hN�
9�H^�{�2*������G~��~��Z�w~�k<~棨K ^�*�^�eW9pPQ5$��D i).�	�ճ��Ĭ���-�^���\Ö�j�6�z|'bע-WW�E����K�ľ
��gAL4`�Ơ�6;}��R*�U^���j-mt��8�����Äc����TY��8���i�ZѕȢ���)�'"�5�������eh�YhP"����c4�����˦����� D��]K�e9k^)՚v;��?�j/`�64i�|�[kQ��N.	Z���=WRȣ�I]��I��v�D�*_+���!���-6�0�ֱF۲n���ѐ���C[�("Z"��)�A�H�@{3�c�� ��ԯRA,�@X`uXҟ���8so�g�����#I�ET�;Qev+ZY
qҾ���~��v�O� �=��G��חiG����پ�6[��s�\ ����}���mv���֛PN�ҙ�zbٞx�u�?n��8
E��Q���k`$R6j�k"���������"���A@|������2�����0UʗJ����VB�>�iw��I��1����횫�(ȋ'�X���~x�>S�����V�BA�{�"Lw��X6d�N~��u��ڏ���n���+���_�`��'쾇O؅)7kk�o_��9{��-o�������7�Ͽ��=yt�jќm�'�B��r����r:q���ٗ�a7�p�]=?��ʵr�^~�5{쩗y���[�B�U�-�'>zB���v����x�^>�HF�ж���j�me��גѽ;j���ߦ��m4�.�$?<9�w��UnA�:8S�LA��$��#���8|A�iv�З����1��k��s��mEOB���и|�;�v����.�N*�*$�	�#_��[@Iށ6ЙVMC:��}�	d-���P��}�ʶ(��N�5�	�m����V�G���縅�L���$HŶ��Q ��Vz�kЮVm;��#�Q�@����䖤��a���V^
�V�g�xYE�f�ߋG�c b�/%�g���lcc�Cja��Ch;�uD�[J�_)�^�Y:V~Zm�RL)�m��o[����X�:�H����#,Knp�/u%wP�>jL�<�P�5�|Fy�M��z���mbb��Dj�Z�r_}h��y묥�_�ԧ>����!�z�U_qV�Z�I�
�r+O���t~�5)�ؔ���,&�g�?�B�ȹ��'�a��%� ~�<|9.�)������
~ %1Z�z�����ҧ�}a=(.PA !�&���#�4�dI���s�YՇR�9߫�a>�2�:[-y��M���k�����^kfúȗ.��zjŘYSy�,	n	��ݥ<�K ����G�ټ#?"��DA�sO���@1ہ]�򒾏9��i��Vf"Ϊ�υ6�"?���t��0�UJ��RpԹ!IЛ���*C��<+�b�c��Vz;@�Nq/���v-���V�a���
mڅ�t+��{l"m��~�M�E|NR��eů@�5Ebۛ�lv2j�>f�^����i���=��Y;x�{�ێx ji��K�������,D�O#�4�O���(Yh���)Ӈq�y�G|Q�눝[�ڟ}�!,2����2c��*L��]B*�ȤVe	�X&�Dy�⊽~f�n��ZK��Nc����n�H\*�,z�c��`���pa��g�X{�<�/J�@��/��})������`x���l���������?bϿ^���5f�)�M�
�����=�ȓ�8B�;/��Ǟ?e/�X���x��q[�\��={��o��p�쩗����=o����>4�D�W�1��9X+���̢���'����m�y��h���[ޱ���$B������L�.�z)�r↋a�{h�>h��Nv�rF��(�"�ߤ�� 6)���*��.��&��Oމ1.�!A���wpW��
��7�(]ZV/����Y��L��P�vċ�h+@Ǝ��A(y�Dx���3%��W9b']t�;�����+�k���}�S�?��������9^J���V{�\tj�$J}�i�	����1�l�*J��гp�J�������������Q��I؈����;��͏i���{X?8[sE_
G�k�1�������,>ˡ���ʺ�[����Dz�Nȟ��@���%j�:��@xhŹ�i:+�ϛ6,�ݑ{���v���Sv�S��h�o�ڧ>B���'/�b3�[���|�2��X$�� ��ȑ�R�v7�i�3�Ï�x}�7z����C����=��~�7SG!V`*:�<H��o޹�TzW�\K���Η
�����*�E���g�|%����r�ף{o~�q�؅�{!��w���NDAY~�����R�Z�CtM�[m�ZJ�$�$T�;�=������{o��`��U�?>S�^������L}��,�j��f}�flb�lii�&'��~6m��;�P��������L)a[��ɞy�U���C���#d�޴���^����m�~�r�>T]�ٰtH�����>p�����j��9{酧`�a{�;o��Y.D��d�'_���
Z�4J�ĭk���b�'�����{��V�U,�&\�����(yh�Z���������v��u�Yj�k'Nb��yG��8E;.�E��sg�b��������ڝ��0�Bv�ܖ}�����x�Nc�E3S0��%��>�jv��sv�-�Pzv��,�6V�ʔE�"G��U�����k|��M�Yٲ'�=n��x��r�~�ny�_s�=���v��lv:e?�S����l|�oaڄ����n���0�Y t�@�j�Ʒ�A0�JQ��)�����Ѿ��4
�B�q@x�pH�M���7��D�
�e���}�5�$�ťԊv��FX4"�p�����CA,dQIq�;r(��H�Rt��/\��Q� ʠ�?��!�W�ΐ��Ǧ�񍏆q_uB6P�>�(H�V�u������!h�����P���axB�T���qc��(*�I;��#� �S��o)Sp�����"��B��-K��G�����5r���8?�Ne�g*G���s�vR�� ש>�[ׂ�\U4¨vx`2PLM�����4d�}���Ox�]V��Q��y2���e��z��X�#�읷NZ����o  �`�=�d �r.���H$��Cc\����+�%�����+Ic�~kx����G(��F��ͰA{���	:��B4/����Ϻ�9�ǻ:_9��z\���a^:Ӌ��[> jp�]�Ȓ��*�e��w��F�{th���9���ɪ�{���ư�Sp�����#��Y�T���!�vX`��:��{!����d����ZJ����r@9Bl�߰��]!R_)}b뾴vi�b Z���me���?�hW]3�LD���&M� &�1���>�����j�a��۟~�!�f���{�["�jWsvm;}��]\Y� �{�6���O|�N���ͮ��h����<�>�w�y����:Vީ�Ͽh+W�����J��5��.�5���?�n��G��뮛��+�v��E�a�&M����J̎Y��J;5�K�O���m�6��j��u[��6�&��U�,�잛��~��v�UX�mR2��×�����?�����,;>�����(p�7:���͟����O�b79d9���f�Ν�Dp���۾q:g��?�}v�Ӕ�1�m�>}�N^ض���"��#!���bm��<o�����g?�~)�E1`vz�i��g�ճe�NĒB뇡���@8 <^A�F,�x��C#@И�9%P�
�p.0eQy�#��=��(/]{�"����)��e]8�:^k�_�ʋ��=��k�@"�u� �C�:������xرb)S�T��]�W�#2y[5$�S�6�ٟc����~kXO������S�+kXק>�H��`�>����O��[G_��<8|!�Q8D�x��<�4Jߊ�hh��zś|4�C��p����;Ia�;���x oߕvJP�?U�F{�$x��ӿ��C�r�w�O$���䗨��.�(�y
�h����Z�j�^k�n�jo�R��E~��~��b�g�ц�:n[͸����8�-� Ɵ���tE��L�j�Q���r�C���4n����o��G�;��tV���^s��E0*Gwu}��ۀh�~��>|�߀�C�#x6d�{�	��}���=��w D \�^�?�{ܻ|����Էh�p�V{@|��D�zWC���ޓ�����i�~����
� ��{^�ѷA�B������nCr˝{�����J}�2hޅbֲ0S�j�_����ʮ=<a�  ��v�w���?��]��[*S�[n����" D�=9���W�S����[n��������e0]�LD��^�sgW�C���9KsO�K�3V��gi�W�E�e���%��}7�q��c�Ҵ�X�渵9k��a�A�ص�-�����ʂ� ��hۑX�^��O�<�E?�x��c�D����%�{?�}v�B��p�l�Gs����g_��v�º%3ڒ>%�L�f�e$"�#?p�͎cU����Ë6?�h�������O&����>��[-��Ȩ	==��y��c���V���,����o4���e�^�h���w�[n��k��e��X�������c�0�)h���K{���4"��%�E���E��3I���s�����Aj�x7z��h_ς-�$ЄS�����Āc�:xOp��d���,�=��p�����B�PBH���A1g��<u����|ՓC�|�L`�m�0�p]�����w��ꡳÄ{�Aԏ��r�;����H�����,=��)X�]�E9q�$Xs���E����辄��I9��,�(p�����ix;U��>�8</�q���D�*�g�����=e��E��i����?�h�����Y�Ըl�]wh��yۄ%�M���o�ڧ��Sk{��m�����ֶ]E�B��� �������Iab�@�|���P ����ttg���=���X��Cς#`�����C�p���+kΞ8��oT���:��A�d�
�Q=�-����*���u���Sg]���z�{J{��N"�7��:�L~\������0�a]uvW�y��/a(� �\��zo�'}`�����p�p���G�\��~6j��{~>�4u�3D"_�H�Ν?k�N����;�̗tK��.�
G&�v�ҳ�%���_�g��[n���l�Z��G󓿨b��� �	�]o����������>p����`{h)8LB\^�ڟ}��v�®����tÒ�\�|١�);tp��y����?|���-G�mw\m��<�=���v���i?�\a�8�*��X&c;�-[[]��{6=��r�Yn,a����>����1�e�S�k���~�F��p�ƒ(�]�����Wl߾y{Ͻ��^���v#m�j�J���w��j,���?K�������k��~����{���y�LʪZm
�9�ݰ���C���]K��3�]\-!��67�s%B!�X���\Q��tW�������׭��Hz֪XZ��ܺ���P0q1_	�`�Gh0J.i�<�K���}�i.�q|vG���P^>��
7����k�I�ǒ���1����Y��u8>z����U?�zz��]�4ŵ�6Om�]��o���S���D�r�5$_g��y�@�P<��μ�����O����ꦲ��5E�ZʵL���m�w�
?`�\S�^�է�j(X>�RtS�ǀz�~�C�j*_�0�^��R�%]�3�U�<�#
�6pU=���S�ς�����n(Z��.��Vm:�|g���|�v$��^wx��v�x0����O>��G����/��M^vz��������4Mz���	i��/�q����p	;5A@����B�����e�:����^�;���#@��&L�z�
��gW������$��U�\9�5*[��f����{���=�?�������+���9����p�{OA_be��\�򸿔ꨃ{�����D��
�Zt����p��#� ([G ��Oj�����/�u\��>g��@��tޠn{ᦌU���wp�Qv�%y�����w�k1ܠO���Q���FzeP��Sx���I��|�6�0f��y$�lV;H@X�R<����ۿ��ۓX��~k��Z���V��W^��}�,D:0m
:VL��Xڲ��)L�ꐀ����=�������u���e�cs��09��BZ��#�LN���a3X��1:�m�R�g_�d�=t�v*�م�ƴ2Q0A�s��lq�����g�6��׆�gg�T5{�Q�E���S�x��{���jm�t�0؈���%��#v�����qX�	~ﳛn��^?[��+k����,h�ưk,C;�������-���c6^Ԃz��l������#GmP܇��Z�޳��m��n����O��%p�����k��G_yھ���S�[��h�����h����Jz�$>���3 ��@��
�B�7��������)��cGc���xO�Ώx>�'+��Wy�{
�6T�/�%C-d�U!�#ț���>t��o���<G���lT�����=��g�M��~�O���|��%��5|O�1A�.\�͞:(�����࿰�^��U>�>��>�Uv��S�)����d�z�{�'�u��EK�h��bX_���|�`S������o���j�4dJ��^o����P9�G�*_~�
5� (��E����lm���ڃ�v
b"���'���Ok���KU{�s��AC��X�ձ6ڝ�ớS�@s�P��u
����!�a-\��+4���o�\��G$>5�!waƵ�螢j83Tg�;2c��~_ ��Y@S]�i�7������ʷ~�mp��Kp�7A���e��^�ˇ�J�F����}u.�x��e=p���p�tt�$��!��Dڵ�����3BC��G�57�Hr��!����Em�Q�5�~tP������kE��A�F}���h����o���C�뇿a#`]��� p�o�;�Rqm2�����L.,�1�>3��նg_�ٿ�����6J.Zt F���[��Mgmn2���k_QFQ�s�6���̅�����+��󫖝8���&V�2�/a�
R<4Y�?-����4�Sj�}�/���o>cw4���j\��&�0QE:~�|�Փ��c�^��"����̎=�K䝌w�]o��n�
����"i��f44�#�=�3�ץ�T�S�Ve`�?{�.�����픶l2���B�~��I�B�BD�M=�V���~�>��ǭi��&����`���v��V}`I���XE�.��?��7����r+a��}M�Y�)/�����
.�t��:�p�iD됁��;������q�C�\G��8(/����kS�7L=�����(�qvx�F%l����C��i�|Gt�{��w�g:����׍3�G6��5<��K�Z~��<L�Ȼ�^�It�yV�/�?�F���s(����	"A}uʄ+<�|�v(���A7�P��:�1lcp�6�`�����S=�O��b�^cn��4�F鼧B�a�c�V/��N�*;�wl�\��n�2�[���Z?i_zr�~�O���k��Z�*%9�v��>i��%��^%5����x%	1/��' �Jh�t���L�$GI �Ci���'A�4zS��<����]Iz�ʻn�������<?�a��÷�q��a����T��s�{_GvN�^W��5|�5��*vϧ{��%�)d ��9�z��I�IA��r�4�G�|\_�ZC&��<�8��f������5e�$�H�3RQzCO���M��N����ɴ5*e�`�d����mЩ�G��ȁ"�f;��v��r����Mv�U���ǧǭ�ڵ��Y{�]��}��6��n��V��斦-�������7_�/~���I���r`V�Nm�-��G?p�͏���a�´�N�,���.��kߕ�ѧ^�Ǟ>f�ܵ�݌V^j�C,�2���f�S3kVm:Ӵxߝv享��Sk��=h�U�u��R����vڎ��mj<o�<�@�X��&Ө��nЇ�4e���բ���?f�٧,;~���Z�v�~�o�O~�n;4� Nf��5��&�-����s��o��u����A����aG��I+�oxP����m6=���v��c�v��/[5��D~�B�]��L����� �}�y9�(Kx ���ܻL/{���w�V9�e.�p�v{����3'�b�Gi/��!����8���ʢ��v|WT?��a^24�}���2Ft6Z<(���|�׆b�;� E
v�ʾ�'/a�Sps��z�πEP
iO�}~Mڢ7�(���ò4O���\�0�@���mV������Vq�ϥ���M.8�,/�۰ݍMK�w��ۧ�o��ն���}�5(��e	�?{��֊֊N[�շz���L�@Z�OD?�d ����]aa2uGUuЩ����3}s�t���3���Z�]p!�r/3�����p��F���j��']��oH��
��rtO_\n���P�(]y��7�;lÞ۞k���Iڛו��T�=�}9� �P �M���'�KI��'�V�j��/�����)b�_C8�Z]�3�S=��#Z�b�Z���k���Yk`��-��P��N�n�xߺ�uk(�m.em�8�= 1d�nP2١S�TZ��0,�H�j�N�ƓX���U���2;7k�a�! �};q|�z-Y��v,c=4I7�7��W߰l�����B�x�P��i�k��Ǝ�m��h��B����.�r��3��H�BSe�F�)&l��a}tB��O��֮%&&�������ҊM�����Ŵ�̌[����V��M�M[(�ME�uQ�6=�EF�]��zҦf��s�pݒְ����X�k׶��|�j�ܳ��9��Z\�U���-�~
n��zm��4�l*ڦ�����Ĵ��3������(��/�Cǉb�	��KF$ghN�������uO
�<��^����I1����%��-=9�	���J{��^I8?J���F���їΪ��+�m���R�u����ABq"�J�ɟ���o�<:�ʦ�.4�L�r�M���ӻ�-��<�	�������7���e�%���衆���X�0�[���� ��a��'�AK�����o��E+�<b�kw�P�_���l_f���b�޿E��oN�n'g�q�	�V=�Y�Q�	���{O�����בp�{���{�;F�w��;|6�N�a�o��%u�:ʾl��%~s�����h9P�e��މ����n c������O��k�;8x�)���E^A�Wۃ�$q���}�|��O��+���j焠��� �PiO}���崗P�a��ڋO���lR�f��?s�h����oPm�/dwً�$�x���1?�3�@ɺ�xX��D�)b�6Z۠n�Bƣ��E��y�*(LRl��2�A	�K`��w��a/���|"�8Vp�r��Gq'+�䀀J�XNe���o������*��ǢM&��H-ԻC[�����_�����4��Z�Y�,��Sf�ۛ���殶�JҎ�����W�+hr!#��Z���mR_!t!8	ni��XҢ���G"�B=��tv�v���'�,AE�c�u�-�TK4����S"���8֙�c��ݾv�����"�0`V<Ϟ������,-(lS�W!�s�o���$�7
�B�Y?I�*0��菾^#!���B*�� w�6ބ7n�G�Iϕ�3`���(����t�Y[9�_	hQς2e�	6>�ܓ��+3��ȅ���ߨ^��k�Qg�U���2��7J�CT
hF�i�1�ÏJ#!��b�*0��GMI��Г>�-!�|M�|p>�^����o|���-��5$�����'��S��s�"�&<#��#�6>X�_y�]�@�+�QoK6�E���J
���G�B�͆+v���������f�9(�[~�M�g�}���K�q��D;�`�@���!.V�x�`lXA�%;���v;W��g��\s����θP@�Bh�t5[�{0P�:](�����Ƈ_��ц�J#���rQy��PH�p4Է7�U� ����jF�D��f���h'�S��+IHL��" J��e:���(��6�U�~w��Z�������`�$��U;_�4D O����iH�� �����0	ق����2h�'���N\������7�Lo=���z�ߕ?g=�f^0=!s�wzA�. $���9/I� q����4��7=_*��(o�-��e��OJ��E�m��T�������|Ջ�ࢷm�,p��0����V�)����������.\��
���Ha�<���S���< �?S�H���p�RRK��)�FT����7�KUA���i?3/�����5C�0�p���-o�=���)Wк��v������T�O���']�R�e�V�}�"'����Ym�'��ջJ#�,� u氾��S��h��V��y��N�������?pfW���r}��=����Hi3�?\x�'�F+����B�Hy�8]����ʕ��?s�Yg�Q�y�zE������v�Q��Ķ�� um��8�
U�Yi����*��/w4����5����Ĩ:����ׅ o�d����v^�CmX���;J��T8,��$�~��hzҷ,�ݓ��[��}�F�
c�5ڍA���]��_��n�Z�	���>�//�$&���4,�{��jo���?�j5�7�C֌�L��?=�F�E��K�&�|�B/�6��i��;��j�PM�rc��\��rG�����pޘFsJ��P��ҷ��� `(���WT���W�ױ�I�<��9����d�y�	���[�+�.�ڛB�Jf�K�	��H���)�%�ȀD��I��uѻ�۞�=�V=�ѕ<<q_)������,�w����1�lςzzا�m��5c	/=�ڗ �D�#�+�ЊS���(?5~4䣚.0<� ��%Du=�lŴU_ŧ��'�U�V.zAy�o��V�:�����K�k}�9��[+Ci�z�L����{�h��+P򆙒[ϒX��b� )�܇I`����?ʚw�C��')��e�����xC��Q��-�+?)�/'tѭ��/���7�#8��r@����F
���>8���W�X͟*��;����#�C{\z_s��1��x��'�+��)�S�r-RR|ޮ���x}�� iqyR��=�Qi�&��I�/ݏ��}E��<�"���L<������a��v�&P<��[�'y(��TmP+EH>�r�W�0	��Kh�/�^�-k|��vӛ�/�r����x}#>HW�҆�R�4b#�U�箔�;���%���?H◺�O���i�@K��U͖��g�'��q+�f�6e���7�L���+��rמ<�lz��v��f4��_����SD +d�8����F�U0N,�`�����Uㅸ��7�;����!iP�6*f�m�PY\��hb���3�:E��u������V�N���Ckn��0B����{oA��x

�l�)��х��"v%!O0A>��ߥ�t�SHpߋ�up�N��#�ڲ꡷���)X��x�u�������y�������#\��bI��\.e��I w
U�BĠAގ *��l�˵�>���!���}�Y��t����٨<%	�C���3��r��ö˚�p���-)c�"X}�q����C�������臎m���^�9�\y��K�%���uG�u���IH�~r%�]`E�m��ѱk�{��尝�SF��"�y�`��U����=�U�a?���.F��j��q�{:+Y��{X��t˅���h���]�h��r���������-Y�o�u�
�~^�t�tCo�-A#����+lYB!��O��mxe����;�Ӯ�7����%9~ghW��D�ި.��E����n�а�<�%�V��B8�U~�+�o���_�O*��#(E�K�o	/.G�����;37|��t2��)"
�����__u}/�}y��s%������;�*(��io�d2�F`@I��
��y� �V��H�}'d����X�^\è����O� �5��=����$�~�6��U��*�흦�ݨ���]��ȡ� i���H;5�*���ًv��y�U�Z��wJdD�cZ�Ma�{UT�d*K[o�:���Wp�șQ�P�Ja+G�$� �B
�]�s!a�����3�k�G@w��?���7��h@s׷��'bm�^d� )�XF@)@�7��_�}C<b�AR��cO�����C�Ο��|�H5B�bGp=L ���ӣ7τ3�Y)��~u%)/}�7��G����7�밦0�a=��@k.@X���J�[N���tȡ6`�A�.�'+��ѻ<	��4D���kٜ=�!$<$8TvW4�"�����g�������Ƶ�1��]���0&�S1�r�h�r�hj��	g5��ʊ�Q�3��`;��p�Z���&V4|<L��k�Q0��;������)�Ñ%�ߢ3���Աݐ��^�;��u�7�A��Z���I�g-��x�$��a>ɢ�����x�Fm�r$keX������o~�C���W��گGb�����˷����k�ppI_E㎎z�?=��+����t�l�*�M����Q�?��"���-�\`���=�f���$��p6�}����dm���u�Y�<��Ä�����˟	�M�j����nc�Gy=KD��Ьڵ:Qk��Ցp�Qy�@�������&��j����5�s�#Cio^����W-�����j�w��}	�`�L�+�ⱶ��Y9������D�����[1
*��m�����T9�ڨ�t۵�U!�Z�"�!�x{�0G��'#�a}k�VV���Xq�'s��zh��tVGI����4m��
	��U1�YK�C Z0XT�(P@
�����0K�ب@�Vw����ZP���f��#�S)�6l�yw(8�ZfJ*˵XIہ����40�H[U~ڏIi�I��zg;v��ZE���"|Gb����3�!��a�Rb�������#&��H2���$�*��������uo�q$E�[���Ȳ���^p7\�7����Į��e��#��U3�9uOw�T�Y����	�aT�4��j)t�.�A�i�q�H?��FPB5L>5����G�H�]
��s*r�)�޼e��[�v��亹�HW��q�ZyԌJ��$�e��3��Y���5�%h2t}G|=�
�|���4*Ωq6lgr:�5G�@Χ����1��0Px�rrM08�4�����W�|�)�^�`�.�:��6���J���֓���v�Q���(����;'������*O����sk�z�Fa��&�N$�MnlX<`���1��9Js=I
�4����|��8Gݒo�j�|��M���r�EK�|�z���d�x��ZŦ�_���o痟�˗/�����.|?��>h�-�܀�fTؑ��9�[7�����ʥm)��;�?��o��!��Q����v��w6ō�]��=%��^/W)����O?�-���������t��pN�E��~h�9�u��˷GX�����C��]�o�n�tO�W����q���V	�w�j;�G鈽_�������w˿�������rp����??��|�o�@��VYmJ��42��w���(�D�W���
�²|���GD�":��^B�aUi�!��W=�x˅]�j�pc &<�3�={��8[�Y�\j%�@��&ja2ܫ ��.�"~�L��9;]�������w6��n��j}�lr����p�Q�����=O��m�[��)�{��X��`��3o��W��񾼼l������j[��u±�A��B�@�k8
_)�F�9�6?h���w�����	��O^c�Z9�|�A��������oߗ���u��P=�g{\�9	>�����O��(��gtcKOЎ����6ւ�������d��p���՝GE�4�堣�t���FF�.�l���9?��Fx������V�2����W�'�<�����U7\[�m���W��?UE�8��Q-�e�������UG��Wzt�|�Б.M�H��@+ct`�Ï?�XGu��׳��w�W�˒���� �Uye�_�sR'���أ<�j9�ͦ�!)���+Tb�#"x�v�싖���<N�3��û7����:{C�s���K��{o�����	��[����rq"`~ZNϏcX�H ���µ��{��ն^D	-`q~~q^����N�=�{�zo�;������h�����!Fsv��J�� ����c�my�a`A��8���-)�1���r�%6�������W��ݣ�>z����W�L�K�+;�XD#���|;W��t��wC�9���q��Sd��δ/���F�\��Zņ$GZu�\6��:V�%jK:�n,W���V������7�?����.��r�Ġx�ǐ�Ր��4�RO�a�iN0���^ƁrN�k-PN�5�(����[��k��Z{����9&A�� o�g%�>�-��1Eo���4���*ܒ\�9G�?��=��(��]�>C��/ �Zhн�P!�����V�pR~LN�լKY�;כF�4�)�ϴ��S�u�)
��t=���=�����~';G
"��Ú�j(*�V�]�J��}�1�0+���R��W�x(\�����=�	�f8
xI�n&{��[�»a �����(A���������_8�W�0u�5�������u|� \����5<2Q�� ~x���.�Fg�pN�D��S�`�L܃kcӸ�
�9t�&���:��8{#�V�:ԍ��ƞ�<���n$��I[�u��D�{�E�S๼8'����4����'��ɿEP�4�3@+��9X#��)e���̶1�m�4-w���Æ��x0t���M���#?M��2`��0ΆO�q���8�G�z��p��������Ϫ���
�W���7��W����ױ��I٘�;<���X�/���b��a[��Ü|<_/o�G�r���.���s{�݆���j���M�FRBٷ|�eA!:̵W�X�u�+��+�rӎ�G��e@
W���GN药kD�]z�F%�.�:+
:��6_����6�Zä�_|����uzt��������߾��mh�y����(ǲH�������,��Q/n+�/g�t\����l��S�����J��a�(I8����Ï!40��	�Dq=6���p
Ùq6��9/�
��=L�6t*L�Y�pD�Ũ�9g���!�r���g�9���\�Bd?K�Zv�{pu5��!��  e�n�?j���5�+A�Kh�1Nw��fo�"v#�1�D��ǰ*C�cpf�RJ�c(%��\�B��kt���H�a�-kr���l,����.޽g�k�p4:x�t����C����ə��?�Rx�c�Ç�و���O��K/����r�
���|�/�KGR�!Mz����������v���E�� �e(/�4;�\#���ўs�z�z�ٓS����� ܙ�t�#��D��u��42�	���流"@�����D���������ot	���Dp�ʄO�Ϊ�/��)ܕ��|��K_�{��f�ҹV��'g�����������h���5-���up�_��r��R����\����҃!w�\'P\ř�_A$�TO/����|�W��w��8��,�?��=h/ޅ,^�u]K��˗�O�Y����n����}
�ۃ�ʡ����cNo�4�����7E��@��δWX�n ��U�  ��R�����%D��ˌ�I��e�Q��D���{��e��)'zZ��b����t9�󯶗�:��E�y���j�E���y�W�D@�����\�4~�\~�B�}%�˰H<�-��6sx\Ɵ�0������lF3x��C"�N�p�ï�_�A���+��@9F��9�A�_G�&���I�=o����)�k{�fs����Z�ş�C)�m �ߠ��QJ_�/�d�`R*S�Rn��B?���ãt���Pt�߭\�B�����J��$b���IW�����Z�_eT��\2�Qs:�_�{�JQ��9�����iTU��Kڃ���sCF���[����p��WG2t��9gl�C������nr�rw@#R����|R�z��'?K?�c��5�q�'�COZ)(娥�T�O�&M��K�'ݾ�2rð U>��h�|SfUӸW�xɧ�S��"7rDk~�Ы\x�OOԉ��E�E�J�ۥ�~�Ssw�(mQ�CKU���v�����]�4�������sD��@��
t��+�3����N2��z���9��e��^r��{=��E����!aKI�g�X ��%�	�&�iM ��yȩ�J�5�W���L�{8�i�=�e�܃ҩ�}o���`�6|��Ͽ�w{�����]�k�s4����m/���iV5l%��F} x�s����(Pt�:���y��m�+�Z���P�6�М4�tzc��F���J #�L������9N'���=����>��+~��� `hpY���఺�OEYAz&޻�/���S�i|]Ҏ���q_�x}��(醿}m�pr/2� �&r&��=C�pU7?ID�ͮ1'?�mcC��%P�oe{Oh�{DC�������$�^�Ó��DPa�zJtCӥ�(N��XX2	o���h�NY���W#P�s��������GҀ���� ���ZC2YY���I�V��%����a$:R�.�[_Y�W�{y8«&���_��(���8�"�9�1�9���5�[����P"���F�tz�d`�(���3��ړv��ϧ�%�@�M��u�-	��W �=ݫ����e4DO��٩����=�ӎ��Bפ��7>f�{�=a��'�ï���ԑ&yO7�7���Җsƾ��+��M�6�q�I�*�H�.�i��,���侪���`��0���s��3杴Ͼ�ݽj�C��Γ/=��������C*��J�-�ٛu.!��>>�%;(!������O��ɞ���/x%->N�#.����o����Y�j��1�7���Ф9^��.-�����^���8ۢ�aų�Y���_==$�0u�|Y���e��r~w�>W_������Eœ?�_��W��mt]�_�]SG��tr�\)��4��K�I��Z����,���    IEND�B`�PK   Y\"U8��Q�  > /   images/86525bf4-9941-42eb-811d-381dc5200b1d.jpg�eT\϶��$Xp��!x���Cp��@�5���Np��B��n�u_��l�������x�ev�=עV�j֪�sV��B�A,Oed$$$��� ���e�l���2� �# ����o���{�� q���'$����z�G �oe�G;� ��;���6 ��R����y�y�y���Ttl-�<]iլ�ܜhe,lܜ\h��8�8�����9�x�����x�xxD��E�xh��Ex�D��  =�Y	e,�?u�����(\< �/=�_�Ϳ2��O�j�C�� � � ����l�GX�W�ߞ�t$�����/� ��t /��z:����g"�H���/�����M���?���4����Ǐ�`bcabb���R��PS�SR��s0�>g���ddf�����a��������Ǐcab�bc��<�|��,�� �#��}��@�CB�CBt4��DC�����QP��1=~�y_����((Ȩ(hh���"���@�C��-�N�n��ܙ�'(��#����DoF��yߺ?~BLBJF��������_@PHXD�������������������;+k[W7wO/o���a?�G�'$&%�|�������_PXT\U]S[W������������kl|brj��tyeum}csk{�������vu��]����v��ۅ������]HȞ�CE{ƍ�/��a�L�'��˸o���x��u}BLϷ�p��i��fX��#��iؿ�X(�� �T����+�G���t������B��5}&c`:m$���=���/�u
�|�zP4�@�*��Ԩ�p;����A�CŜ M��b�1gDK���L� +V�a�v���d���[=�b�c�"���&5������b�+8`P�p��� ȕs��{W@����-/P���̭���p������S��͸I�`b��;ތWL����Eb�&g��F���x�+j��g�(.�1�e$:߉s��_��ջkc�;�*�����V����m�0�z/��W\_ڄ~֡f8%��]��^]w���c�|��-���&�ZH�:k�ޙ��2;���E^��l����j�s���" ǝrB���"P����7�tǦM<4�;�8�wyՐr��[�'V�Is	��!3�T�ޘOs^	���bH.�4q�7]l~�m����}��W��l�+&�VpFhM��E[�4zV�olz�RL�c~�d2<��b3L�Z`8�x�Z��xi��
�����Lox��L�/��h�G=&Ώc����7�u�և74��W�"�2f�SrM�Q�<�����.��ձJ�wE�{c^o�%�E	;�S.�&�Z7��2�:���tB:�-�U���kZD���<�rp6_��eU�/N������M! b8��1���?�R����ԑ�H(s� ���i��]��<q��tS���V4��:ܻ®퍬(��]y�ڲ)�d����"�	e�*�0��k��ޑ�U�.�:Rv�1."�l��2|:_lID�ғ����UW�U[n@N�|`{�󧊋-|�����p����wu�����=����H�ٿ�H&ٛ �\�[�0�ڋ�On���d���ɼ:=
+�|m\Y���Nc|�u�������G�����7
9J�f�B���Q'e��Vsq��X�e1�K}���dzQȷ������ҏ9�E�r	YWWa&���7^/�D��3�B�0�)?�'��7u�4w��7��ֱu�m�|��ý�36�����hZ����BM������{&	R�ㄭH�p�'��g��;�CS��H��2,����D����F��1s�M�tG9����d�a�"��m�X�v�Pa���U�5E�������LA�Cmv~���fIO^7�u�
� ���`R(���_���zX<��qEP�|�+����4�3|J���)��{3>,��ߨ�kO%�>ͮzBKW����X�WT���7��A8ۏ���ɡ}Ы~o�eŧ�H��#a�m�	r������eN�(��/�e��.��Uk}��rK۪O�(b���78S �jᰊn��H�w#��/��9�|��l��c���ft�fk+%	+P1}yf��Q���u����_��,u�a\��.���ꕺ��h�B�}���\���4"z�>�H��,�nR	ݞ��b��/�/p� 'G����_u]_����J�c܈��캯�1�è�Vӏ��.�H>|򈗷�\� ����)Ȩ �H�.i
�T��3C�ED�N�_�$X]#�L�]�O���J�6c�Q��G���+�C�y���1���}4���|(�KAr��.c�fg�/e�Hp�g�:MҎ�u�����B�~I�!L�ǫ�)��٩��i���iP3��F �޷Q���d���9���f��
��g�ꟃ_�����r�o�|߮��h��*Vŵ))6V�4���;�%��fˈ�k�M�C3�����"&�Ye*o$rO�i�D=]��7�yO@�$�c�A���9���Ua�|�A�)1N���K�%2���5��P�iZXĠV��5�D)%�[�N��l�s[حLq���h�?���|T���������k� q���Q� +���A��A��~���iIt|.x�y5�	ho�A�-#�Z~�N�)8
��J�yn�Mp�i��?%�2O�F�P%M���Š�>̇t�J|4�I%!7������Ŀ��5��V�4���_(E�d�� ��5 ����>O��kl�&?�|t`+���%y�S��i�?�%15��/%o�ʀK�>��\%\\\�A�_��z��t,��,�n�����6��v�����?�XRT�oEBw^n��zv5��xW���a�a��5�����~Z�8����1_'�K��׋�'�ğ-}�~l~s�z���C�v�&吧��$:��Vx��*���F��c��-�9]T�w���N߲,�|�5��(TE�<k��"�:H_;�w%��_�
�]�9��B���G��M���J
w�짘ꔜ|:f������||V�����p?�s���l�o�߾p���9�D[���/)1�K�7}��O�A�D��sW�MD+� ���3vխS36]�c�Hq4�C�1�L����q�W��X�4}1�V��KWЏ�8�J�ɋc~w��F�
ΐ�Ds��gHQo�'o��Sz�����GN�Ĭ+q�N
'��)�D#����+�L\i�l+>꡾�*�?AO�uh ��I͟ZkԵ�A�z�GG2��"as�Z��s*�n��������I��8��ANU�pU��Mmw�/���;�㈊���1R'"1��S������*�'� Q�t����?J�.��dY��;��Sp�\�,`��(����1��w�k�p=�~�.���I�Z47�����<"���d�H5��]w�F��of���pv�������~=P*N~#ꑅy���3����?ԧ��v@/Eۗ����;C�SIj��
��mj�� ����ݫ()��a ��[v����~�9^�^e@���R�qnN�N��:�id0S��a)������QU\���iKu(��O/���b�у�Y�3��h��\Z$���a��h��C9�Hwf�&5����'����ȩ$I�BK517Ծ)�S�@�7�|��TR����UX �`��S�gZ_u�i�>F�i|���+�U&N�:F�w2nFb؆�c�@��F��7o�U���}W��>Z/�cMn>������훙�p��$�P�Гf�F2U�h5�Tx��P��1;�s�������Ӥ�'��Ǜ�h������ךeN9��e��.Ndx��E�]?F��Y%��k�`�P��_m�oywa��З���5hX:�b�݀��v�p�\�9Q��>P�U_j�B����aԷ���*�R�-��ʈ?sT�^ں�!�3~�Оp�	0߳.�6�$�K?�c�Ť
�S�x�w��L��l��2gf�B6��v1ݶsE|^����U�
��	��捪����� ~~"+m�w��6/���s|��Q��V�s%��0uM��v4�~f�ٻ�-���V�y��(�b�6i�	�GekOՎB�[�d��֟	E�(����6L.ί�e)cd3}�����l�}=v_�D��tW�3 �Μ��0S^S@ �'��?3�V���S��ƃD��&�'O&Å��D"/�p� QyY,� 2y+y�"J�� �T ��T�[O�je��l;�*�q���w \��n��!�+���x�V'���WV�������k����Z�"��1=꜀O���*$����������k5d9�O�N�5f��u���'�+;�2c+63^���@R���H�a���"sJM�:�����绣N.�{�U�֗k��@�@�s��J��¯�B��t��4��"�3^�?s3ʁا��O5.τ���O���Ϳ��CS6<�� ���-.}��!�u��
��<�6ǋ@�yt����g��%���'�������ĸeļ���<i�D�$��̢+��Y`"la�)��*I͞�U�~��3�1�UW�3:��K1�1t5�ԃ��x��-o�٘;�F���sL-=Y{��/O�z]$j�R�#w���w/|2'��HW��.b_Ȃ�7�H�z.̟+�u�z$�7�Q(lN���
=T;��V�(8����#�fߙ%ցrJm-}��HV�kH��'�����4�A�&T,����e�Q$��D1��+{xz��G�Q|D1�2p����zـv2�b��7��BZ��ɤ[�+��~RX�G�y���>T�u�y���䄪���6��K��{	IB1��n�y{[¤芡)�. w�
P(��,#�K�Sa9���n!�\�������8Ή�8m����ݗ$�k�]�I�(�gSf=ń�,�yh܊�&�@k���9���a��+?��(B�J�a�ƣ��2��fB�~������J6�����I�Jga��݅:���b�왎��7����@�:E�+�r��:؄K�# ? r���1M���DW;���%���PqI�']���j�A"����ܙ��~GmdYC���ňΣtV�<V�f�翲�I胂NO���LCJ�~�K�$)���������f��+s�s��0�}/%	kt��^/2�IQ��c����	��w�d�p���&P�3��37�hjJ�|���G���;L6�u�"�7�v7�J�9=���y�@G1��%�
T�=)U���h����b����s�{)|۶�7$�X�|/�@���ձ��a���ۈc �w��.|H��Δǔ
��R~R��U�¤��9b(��������f��A(a����0,��m}�϶�~?m�H�h�(�$���sZĲ,�T���g�����9��K����#��3�B`}���?���֠��u�{��*ge�lￅ����h���]X�[�D���%��t-@�*�^���ُ���ն�;H�gz�KהӠ��W'��!f4�`N}S_�Li�������� )h����;pJ��>��1N{~�%�Ａ��Ox'2'�ZɎp���E�&�9
$�*��Ȉk��	c�0�7�z�e�ed�S#�������u$o�
�;x;36�|������H٨���w*j�K��x��[��!��53�>�V���x��h�;���j�*JUY�&�=�ׁ�S����JF���b�
��y-���b�[.ۺ(�YXTn	~�����߽�.�9�,Y{��(�\��P�LZ�de�(x��%ɮ�o�J<�-]O��J#n���&,�l}�Θ���.f��ޫ	.����/�x·�h+�� ��/��kْ���j(�\���S����d7RaJ�䤫��2o�-�s'�`��o���o5�9gڍL:! �������=u4u�J��yg�p�OC`��rC�JZda�8_�����%iN,��J��ͼ7X$�|�g��p�,I-L�%(�0Rs�=��7���W�����P�!4i����
	�ٙV�G�q"8�'W,c��:�Ǯ���n��)�K�$}��B<2ޗ���Z|_���VC��"�D2?������q:NUb� �!G��RƳ��f]�NA�ȠaE�,�P���ո��#�0�\�{���U����~(4ڸS�O�lP�5M�F�3�W'S���с�a��z*���A ���'�2\��x�e9�r�	�{�_�<��?kj���pv\3|��`�鄽7+"F.�h��,]�/R����5�@����$ۮ�<$�?oN�P���kF� ^y�ϱ��A�;!�^��������z�`���W��A�U�ȱ��D]f;m=�:i���(���e�Lͯ~���ҷ�-IԢ%�Y�=L���ŜLM���.)�xDL)���^7��z_\��y���2�(h�c�>J3�3ޡf��;�8#8*�z	*Rw�T� o���2�.����*�h��h��i2kS[я��ґ�@����X1��# |m\T�������Y�k/�Mq�T�0f�C}�̻Xf5��I��[&��ʶ�������:����2N1��m�����[aOq�6@�Ք�iC�ށ�� ���ʪ�?
B"S���Y�e?�]�����'}l��6�=�m��C��gz
H4SE�;�/�fOQb�љPDj�DK>�6.׆����[��# E`$���� �f�2o6=�_��	���[�� u �j6R��9�E�����qbaS���;�����d�m�Z��G���V��V�/y����Y�~;��<�L=��v�By,�z>�m6b|<ȯ��6�df������etδ`����jT곞�D󞰨��/A;S
��c`�uCB\���볜:�d�y�缬�dя7g�$){#�7����ud~\\hdڲ��������Β�Yv�oJf�ulJ�Tk]ZM���"�+ލ�u5�w�1QX.Px�C� ?g޽�3���1�]�l�_`v���B�W$�l�����^��e�(�u�SN�b�腬��LC�ږMam{p�[z���H��Y�,� �����T�xYa�M���0v�I_�/�Œ�,7R}=��r�H:&������e�ă=��e�$P�+f
�н�Z�@���MC���l?;$v�M�]Z�271�N�OU�i�'w+�����V���	�ua��Hj޳�C1U[x�؛cj�'+�\HYvƔʢz5��H�7��)cz�J�tG����|7}�b����XܐMIrcf�FՈ��)��_�|2I��BKӐ���fԺI�¢߳K&Z���o��$�x{+� L,�`��mp+H�sF�T`5��j�w�h�+Ո�����z~�j�T/L��i���lf�|�_$�����!uA�~�4?�>����ѯ�����/p0��FI�<��H��aЃ��b��C�1�Bzi˕�S��o^>��^�?��,D'Y��j~Ԛj1r�������$n�" ��w����g�:�2r0ĝ�t+����blfS�>����ZG���x=���������~G�� ����z5��xGP�}��C%ҳ<���g���0O��9�R�g��5vQ���Z��u�l�+���O�[��6jߝ�S6<��R�腔���Sg�ײ&�e�Q 9G��.�������?k"��N8�
�5��3�8�4j�c��h�2�n��pvSw�VgG�.��9>�G��?g�<���i����Ѧ43�@U�܈[U���PK�eK%��@Y�W�x�?�Q�g:%�"5&.x��5ϊ�0�?c�PD������mT���o`��[1sm���*�]]ތ���Ϫݥ��rR3Kr���F��^<���%��4��dOT����
�BȽ�����X6�[�wdw�;ݟ�d.�I�e�)DC��١�/S�K���8��s�w�/ta����鈳��<x���Q�-06¶����z���^6i%q�1M0����m��i��������ט�KB�ٽ�4I���ƫN�rC����/�#���;���t���-�ഌq�㤡�!�J�9.���!?�'ƒ�G\T��{�vW��6n^�P�^��������ķP�^�HO�ײZ�7�ֵ8��d��6�փ��3߯3U�ӝ{	����/,j<��u?��`�����߉O'����䌻x =�7��H)���c�\țƲ4c	�5h3�y�
ε�e_m�#�*(w�?�$<��U/g?�+b���m#�3Q��¿^8�{-��E������dS�=���'c�"���~�����8�r����\p�S0�+-���EU�u6נ�XώY>���;�皀��r������iY�����{�,�;�����O�t��4/}��u�v�Y����_t: }睥���P�?DL����3�5���Pc�
�g�o}�ѐ_�&(���4ܨ,�F㨪�U�]�L�]�Hƥ�h�9��Dc�O �͈���ak�+����Cs�Ѣ���������
��\f�(�5H9�6��3Ǡ��{o�>-7���M׾�>j���z�$�$�<�H��Q;fV��V����,�QTv�#��3�_��S����'Rl.JH��ā�|��G��iJMI|ށaZ�$j�[�]ǅگ�=�y���	z9��Mt���#��I��,K��診�X(��>�HTyp�i�5� I|k~�ە�S)�aAf?��N$�#��G��v#m��gZ��2��zD檂.�=��	4��;��ۂW�u�F�r�\�;�
�yRK������_&�	�Jy|�<��<^�S�iv�d�P��������H�$�_�[;�������3�13w��qk;�����Ċ���U�F-�\�|y�蕋��/�UP����}�dn_�l�gd�ne�B7b���;ݘ��6�3��e�'�R���)ASs|��ehi��~t�եw����;fWV�k��=����v3�g���ّ���j9
%���l��;�>f��,�Y�eY�F�$�ڛ/Hh��190�#��������o����\~����k�	g�\�{4��F�r�����zugwtFcw�z�j�SKu�cH��1m
n��iW��U�{��6B�';�.����H����u�]�'.�45�O�#[uA_�	+������5>q)��ʽ&lH<)t_gل�,j�&̺�a�q�8_sd�F���z1�F�1���.����u:9�uzζpT9n�c�U��;�c��'5o�F�1"o���؏g�
���=+���L���e�3��-�l(�N�����T��Z�|��H+���*9+�>�oL-�Qen
s��F�}�`��K��ty��s�u�m���AU�9<��?*���`�R=X��>C O����(�[uI��B���碱�Z[%tS=~���hKI�b��F���īYG��G�T,����
���c�fr,�ͺ?���8PQ%�lJ�7��>X�qܞͭ�P�����;�s��������ټ���\{�%c��͕����K�B[uh�W	%��P���jz��FYU*�D�V����L؛3K�D�-N�>9�J)w�m�C�Ym��qbdXΩ�&j���Ů��p�(K��
]Euk<V�*�4~s'-���"�X\��MS�e%8�c�����#����m5Ok��� m0�Y��J|��:E��j-��CC� �S��2��3�/k_߻�D�Ϸ�V��GSS�!/�P=�G~�F�Y�  K�9�o\� !�)+�z�]4��-^�F��B�}��A�cbs�k3�����m'z)Т~��y\[4�Ǜ����n.^��G��%�I8	����,w�����{'�r��O5��X�޲vs{/�����af��֒��Ɂ���='7' �zofng�F�����Q�񰹍���B�Q�_�K�������������������#H�������{K73Z/{GW/���]�^��4�s	1�w"o^����������ӓÓ���Ŋ�[XX�����������������+��+xe�j�b����ɑ��c��N�n����m,Dޙ��ka���֌ׂ����̂��݂��B��[������h�����mW���ˈH�X��9�h:9�K��~� ��_/�W=����$���!;�0;��?�b���-��]���8���?s߇��?{���i�?���� y�<@ ���� y�<@ ���� y�<@ ���� y�<@ ���� y�<@ ���� y�<@ ���_�ڰt�g�dI�mGad俞��z�D{��޼hO00�a=���|�������)�S<B""",\RbBR|B"¿�(�r*�c4�Ǆؘ؄�������� =�Q��;
߱���9;�����껛JE$B�7Tݹo�ݭ�C���c�^� ��~��n����g�Sy�uϕ�[&^�	�G}y���_'w٬C� ���r�,~^�0�����*:h&�	�/���G,q8��ң��a�3�T������=��ؙ�W强P7�p����ա��$I�c��m��J�2��:~(��Rݱ�ߊ�\|D ��`Q�H�]����d"����L��6*WX��M3^G�����.�X-�t�s���
���A�:�-e�p)*��=]�,�	a���hj@wD�����)N�t#� Fu���� qA3{<�~�۳ x���g��(oN��f �ٟ�lY =�˾�S�����u�_j	�J_$����Y�F~��,�C ~.�fw<v�wy�|�X��
��tU܂;�
j��$ĭU���_7roy���`v�M���2�qf�T�AAAw2�6ɝ]Ӫ���?'�G4��CuV���'���;J��GM��a��(�h�q[���p=�6D�I6���d��� Λ�eʷ��.U�\�)z��֊(�5R-�x�H~�����Op�|{�~�
O�J�[����=?ޛ�~�]�Ǯ]��h~�'?�� 1��b�9��-�����F�Vw��VF�s��+�W�@y���lI���.�+��������މ���[�u�!��x�@�� !� ���F;`T���& �ؼKG@��'�� �>����m�-�g1/b�5�]9��O��;{{ʥ��O^�x���X�x�^��NU���5���O{�0)m���;�x�y�䪫rwD���E6�fؘD�A��]s�V��_ۅ�"}��×�予�s����ћ�MV�i2�m*,����A
�5t��([��2F��֒��������0 5�1�a�;}
Xl�J�r
1i_��#w?*D��I�wPx�
=�ңױ8����!7�m��kre�&5���Ii����NO�
t�Q4�L�y�^Ӎ ����^�w9�,�s��&]�������4}�e���p�hƖWZ�Io�q�7Vu�痒����bSF<��^�ΐ׊�H��.t�̺�(� ��hjT?=S��X��TV��B�������w�lwt*�Z������� �+�^�6�  �A�[�Njw�Nr?Y��}vZ�`��۩��b��-����W$~J7J~���ݜ>g��6��^����� ӑ�oJ��ն�8��t���r*r��Y�͑iq;%��9hrʹ;�uc9pc�*vۿ�!��g=.�f�{������l#���V�:T���Er�09?��7�V��:x�w/6���X��N�Q���n�����Zz���Ra��)�TH���,�zv�U��tVe�3ȁ���W� +��w��e>K� ZEnt����Ň�j����AFǝ�q�L�73�'��.���:P�h'��R��o�g ��M�9m�a����.���
�����{���S�V�TƊ!���Y�@��W��ȱ '��E4��˔�G2�{9�(���S
�8wIv,�6�����r�J������S��"�8���?��Q�a9/�^E� �x��8���4�L�9n��{��Y:���t\�ّ[^�NОm���⏺�!P\��\f����WL=~�:VJ�7�~��U���n��P�x]=)F n+��_�z������)��V0/8�Y���-��5��y����9^�hIt�o�1V�)�bL�]OrC�,1Ȁ�!��!u���B��C���sP�B�������ی���M'w�*���q��wr�yj�8�BW����J�h`�'��~U<�!��>m��2籂���ou�4��*<�g��sU��=���xd��1�>nBy��v
��V�)�	�>���KF����A�e����=R���G�v^�o�uW��M���op�@Xl�xvC.�4p~���}��-}��VN�Xc���l�W^��»z"��i����Ζ-�2�	���R�fo�s:Ԓ*ݖ.�>!ӟx����*<*J��:E9B�
��l�����?�x~B�z[mNm,�|%��ø�"����k_	g|������^�:��'C:޼�KlO=>P��F���0r��F�=�:6#=La�G�@���9�hF�,J�REe����gl��z?"c�2:�%X�Nu_���F�;%T���^~�c��h~�3?Nۈ *���ؿ��^i)D�`�҅h��t��)K�h
˪�Ui�C A��J�Wq��O5�l��E��=^p��-�
y}�x4&m�ê��3��n" '`��чɩ7�F��: �}H�]3A(�y�n���Ig���=��q:l^��w����R^��W�C���n�p���  c\�e�Y����w���,�}%�ǹc�vTZC�6�d��'&���"���=��G�6��Ϣ$zK(���0�g�ri�N�[Y�~=�������_�H�MTRAHZ�Ic��~�G�{�-���vQ����|��@G�8'�|>�qF6=&�w��n�Y�{r�-M��0H�=��O����_�6˹����c-Nc�D������|-�s�vwDu���������v+����*�r���ً�eX�l�0�;�Ds˥�sC�H��O�ܷ�����%�Uٽ���Azb�Y[�@��}�X�z�~�0JNռ�mBt+�l�K@C r�s����5��N^�P���Jh�e�DKo4;7-H�u	D��=q+�V�N?33'���x��M>�+I0��@��5Z
V�ڈ!�<�l�&�����mɿqx_��U�փ���D����b�?K��O-��X0�>�bvZ.[�'��s�l���/����� ����W1�W�?��&R���(�P\��庉�4�9��y�Y�w����̝</��1��
�2�M)R�и�����^��ꀉ���՗��$F���e~7��w��-�&w�Y��Y����~<��!P�pئ-�"Ǝ_:#r��U!�g^~���Sڅ4�%z�%�n&Gj���d�2��r�7��'_�w��Ƙ�T  �m)��u[-�h�"�����T���l
���e�*h<8�îk�:����&�S���r�TF��
-2��@̅|n���NLT&�D�t��M�S�������)�A�([w��)�w�b�7^�����U��{���* �f�G}zO��{40``�]U����9��0G��ء��<�5n�J���T�;������<w�a���YF�R�Qr�u�0r�g��5��U;�g.l���l��x/g�DV}��J]mf��P��݁����gz����0id��G�E�(W�`�%�+�p�I���7?����xχ3�(�ۅ�O�������І�e{����*\���T���QM�[A �r���F�LF<�XW�@+�{1GU@�"��ËeO��a;��8]����!2U�҇);�K�ɟq�$�}����ʮܔ�zU��F�7�!3a.�o��M~C"�x]�*H�2�[,}_\�>N53����U�વՍ�::99��T�E姮X=���� ��Ϻ�<4�-F$]��ǯ�>�,������2��PZ��K~.�0n-��Ҝ���l}ө�|G^��׉�6�A�xն<ݥ'��3c\���x�E�@���/vEx�{�'*���!�sS�e�D�MZD+�|o4�
0�E�Hl��m������E:ЌN�_~��uH�����MG�J[� Gu�Xz��<�[��{��T����,q�s�+�f���b�UE�4����o\�+��ι�Z|�<ͧ�g^/�X14����Cx�z:
f�B�P�wWlP��ZDO�_�d���7��3ȑE Y�1p����Dg�P��搦E��+�A��"E�H��z��
�y�]\맟$�S.4M�zE4m[������������[,]��F�wWp�is��M98��e��ms�=uL�EE���e~tg�4U��D��X�]�7rf�h4H��?�kۼ����"¡ /�������X ��fc �4ƫ�k�Xp��.`���Ut��g��C�%����P9���<?� 0Mt�kN�Q�����P��������=�y��a�_<����p�$P
�:Ĉ'"���w� ���Ud�%I��~v���ɗJ���tD}���Y)��t�h�xF\� ~&ާħ��hbf�GX�C3x�U�>^���>�ҷMb����'����m�캂KC����-v�װ�P0VyS���f�.�����"ݪ��S({�W�	�������	��o�-^����f���}2��'-e�� 9nR��n{^8]�1�_�ͨa}x�sr��K<�v���Y�I�վ�Y��G�������*�MUM~�� �(Hj�\�?eꏻ4�,&^T��5��ì%$���ۥK^���|Y䰾���R��;$�Ɔ�3J����m�1�{U��
�}&��p�QU�̥��YG7��Y���mT�M�c|�����2�����v]-�o5'r�_X�V����v*v6^\�����@]ĕ��b$��������#��τ�<�s��-�XDF����n!�ٸ�����s�as�@.x�V
>b �4�����a��I1{s�۞��BrN~w�57,/�s����M��mm�^���������fT~;��a���wT�a@t�3�`V�r��r�H�Z1p�
sW
?��T�m�W��GQ���@0|Ȫ�q����bq��-HJ�H�W#�ZNze_�P�w-*[Ϙ��2.*�Z��s��({V�e�x��G:)���S/`b{�m��S��t�77��S>z2Zk��x2^_f��n�o�4��앢��K�ޥ��R�4g�1	���}
KQ���{f�E��^���]c���`}�^�,�'���ә%�k�52Z�n������t��� ��Q�:؊��Z�L�)|�6��Hr�9�%��6�����ZT�{���'K��;���u��$�#ЧE��L�'�����k�o��މ�f²�p����8�x�}�d��^.0�c���i�b��%�&��'o�"��j�s��r&}��*(�t��G�{ �ƭ���FT�,E[]��)��IIu%JH�Jm��c�(=�̎�>I�E�[u"�������'�|��҉��mS���l�u���P;����⌺�����
8�(Ǌ͸V�fl�:�����BFکs�R����%����h�ȭ�J_���e~�Dp�C���$����|�-�Oc�%�w� �Es��;�ի.�1G��k��&���l7�	�Q�$���ѝR���MA�aȝC۝�SǮ�k���D�T_V�UP����*͘d�)<�z��˶������".���&jF%�Gv����܈P$?���k�A��N�ͨC;��Db@ �6���r�n��"�� �����R�NZ�>��.j�o��N\���Z����R��?��2�g����t.v]s�ۈ�J�.�\(����3��^�
��Xq��O=�?���{׍ RϮǌ�rdu]���C-Iya=>4�h��ë���N�Qw?T�����	����S�cN�[��	�Oi�Ie�e&nV���_Ͷ��/7gG�8�)���J5���\>i[���b��(�Q��r�t��Z7��!y�D�߆O�~^���^��g�`F������]�;��|a���1(���v�c�iii{$*�s��*m�B��6z���:��X��4���ļ�������G�g~q�D��b�]�ڸ�W����D�|ߋ
��9���)�W�  ܑTwFY��ֳ��Y�6�DXv|��	��F�p�;���B��D�89�ܑ�D�6�9CD'O3M� �>�5ޣc�=Ѳvw�~��e�:�Gف��[�>r���Jܤr$��A@�.��1�@�8�v��]�����H��g������V�b>F�}vH�K�eǒ� �M�/�)B�~	��3�,I/%�#��)��1�͔>یf'��4}o��&EGt;���do}��8�
w��gՌ��L�O�p��1�n2�1�W�a�`��!8���tȖ�-�~N&8���ƞL���9e�,�p7u���UL���E�ׯ�)P�/�����`�Ƿv���moۮ� L.�� ���
�,�����~"� ��]��r���i��W�ڰ`�	�=�\��ϥ�St1/�$[� 7��$���8� �5�cƻ��3;ml �N�}\tLЙ� ��?�{ʴ(�辮�Z��F�H�Q�QM}ݾ�F@�F��"R���.]�&*�� QA)��4i
ҤK�t��i�k��� $7�s�}�8�q�}?�{%�k�����5g�ځ���?JJնs�-��I.V7��M�e ���_�a�b~(twW2���f1B<9-Y�ϋ���������!$������$q�h�ZxEi�m���uQ�����`Hhy���Vב20#11sU6��#�]������#�dhbU9}b��X=��Y�]��p�W���.w�b���U$�9�\!��W�&�y�>�p6�ʼ����� �h�X.V-���%�~���Q;q�n껙�k�,�����	��2��u�C�/<��$vʧ-���ܱV�y��'���/�tX�:ܤ�d�hF.����wJ�����k���pt���������Lh��R+�e���W��e�ϙ�.W3P�T���^�lL���eIo�$=:/{�l���P�(��Bg*�k�4�F�|����L���k�>k�����k`4@]��GM�� af��ag�)�A���Ű6�W.b�Z/Liߜ��p�ltQ�y���UY^�^⵺��f3a�_$��BTx)^Jò\��&+�i�#"*��!gW,�j;����y������F�B>���̒�g��GiU��J+^��8�noU��0���:s�E�o߇��@��s�e+�2̛�ڔ�����-��{Ω���[����v�
��c��xp�ς
>�T�F{��Yh��ގ�gjnf��_s Z�XZ�������W
�K�����&��]����ת�+v-��'Ģ�[���ē�W�7�̤�.���݈H��a���4E���C��[c�>Ĳ?������Lͻ�6��م?�,����H���5į�4�������t\�ղO�87�e��x��2�n�#f���;h�
wEfk����˩��Yw��/�m��p�&(�ĠC+4��fp���5��-3��~�ToY�@�J+�ȀӠ�>��7.���Е����$ǚh�����*�j��}b��ٙ��I���!XZ�:���ת(���J��}�%�F.���3�ս:��h�p'��wэ��^�+�ZIQ{c�ֶ~�kCb��.��A�'���	BQ� ���~���n��g{��r�O���0��S���Qu�ɟr���.��͍,��]	���+�)�[�m���	�ݼUnϪ΂~���B�
�um�|�\,�q/�:������Po�����\X�!������m����ߚתC;��MG�o3�d:��g��O.��9��譕���B5u�*«�up�puؤEI�s7���sҽ���,���~wɉ���{�W��{񞳽g��	�v-��s��̔m"g�4��kd-�T�K�t�I������L��UQG*�-5�D9[D�H�����o�w���r��N�M_��-�ڂ�ve�Ld�����XU��s�Uؾ��Ǒ�Yh��^L��ｿ%r[�<P�ˌ ��˝��rW0��&W�ј�byw��_��Mu���LJ�ݍ�����aZ�yyXR�.SSV�N�5z�̈́���vθtǰpf�m� ܉�W���ESf�<,�E�Na.�JS����y*��c�g�J��l|��
7'�ѳ�?��-ٗ���g�h���}7m�������ͳ?����խ��tF^�X�Y�p�ք:sܟ�w!Չ�'��6÷����=��^K�:>kS9Z�{e�����hw�Rm��>�����������.�E��,�V���u��(��yL|���M�S���������T����۞?��ׇcq�Qb�����|XL ,�{�i��'��T���O&=�BB`��E}j��̧F;�Q��l��M���t���v+��C���3�˄�e	�����f�zbܮt�z������Va���\[�-=[�c]W��r]}�J#��J����n��VW�#�0�3b*�1p�:�Xho�%���V��]�G6�W��H�ڳwN{Mc!��~����~_�w��cm�z\�=�S���y�a�_ 4̺*i�z܂��	��e��א� k�Q*#����&s ~9#:/�ϔ��Ç�SDk�~��uߛS��]Z	рt����B��kW�ᷔ>�V��g�{��>�b5�c�$���c�����bk�D�^Dk�p�R��f��I-�J�$9��b�7�#�E��f��mwߪ�lcb�~���ӆ���)�2n��59����F;o/[Awrg�Z�����Ѳ��7����W����z���"�vQ�!r�����<��Rpփiݦ ����&ױ�{��y���Ec�WM�/��)��+m5�륮�cZл���T��D�-i2ET�6��+���YX�8o��[����T���1�9ki��vfX��p�-��[�צgX1-�т�Z/�����
%�~������������ ���֯@b�'I޵�o�J� q���d?�!n�y�6ׅ��"��<�xS�Ʒ�Hکv<��83�NW��kI�lJN�=�@Z�!��:�Y?���������=�ZG��W&�(_���*�d��s�e?�}�XX��y��[mPɈ1��������G~���f'_���I-� ��� �&��4��G�d���\���?�Co�Bh��5�_.��a��_���`����1/4�i�ٴI��Zi=�pF:�����7&�X�ɱ�o\��\�����㞬+8�h�it�Iլ�L[��+����γ��z��4�N�ݥ�G�ng�coѺ*�Mƻ�tX�,�zy�v��kh�|��18K�Y@�_v�R'6�
�kt<���A�_��7]��Zi�`�JfS]�v��bֆ�d�גZRJH�;�ܔ8d� �f�O�����>��>8kC^K
���V�p�[�@젅�f�M}�3Z>����m��x�U)��`��r"��[��eo�1#�ɝl5��i��rY���`�h�A������ܷ���r�#3�O"v�`u^��@�4-W�MT�I=���UڣS�)���d���jE���u���?X�����������_�D��g�
�}�����}0P�t8jiJ�3�i�����晹�ts))0�w��tDLPgU�Hm�N��;�lϱ-���11�X�S�}ᄪ����{t��~�ޭkTĴ���[ss.F�e'�xw��w������E��v��Ǔ���\4��8�}�Z7�=�L�/��vDa�VZ����4�]�i�y��cu}s<&/�{�WS�B�]t�=�M�+�	/�@Y�74%�ȸ���W����N<���/�������7,Q oHL_��Y��~a�Mz\C`����m�=H�a��tQ��[LC�|ψ���&��gC�۴��b߁h�)�u}��/Bu�iyr���ޛ�ٌI�N����z���g���;ѷ�ڙ-�)��ȵ�����oLs����C�+zol(ϴ� �wQ3��]jd���ԣ�7�0��r��5�<��6)���s��T�[��h�v,��S_�V�:~E�:�.�i �C�ʆ���lG�K�EY1|Z�.l�U� ��ݫ
����R�;�C`v�C��u���t:m��ЛD�m���Q�؛��M;�h��zOR�S����Yȸ:+�Ij�R�њ�{�HP��@h"��xw�E�9�}8$��31� �	*��5��(S���2����_dy��k�Vr
Iz ��:�Q�:����_,���f^����"y6ߝ�=�wC��*}<���m:CB7��[z�arNM�07d|9�'`9��M�ԃ��6Mu2F��k/7.��u���@��+�bN1�$j�s�;��7�<��?�uڎIm�oaw�c2�oc��ޜEk>���C���`�w���e�r���}4���嗦?�&�{� ��ʚ�oku�ӽ�oiS"��9V S]v���Cf`O0�����R;!��+�/q�I��n@>P	�Q�� ��	ך�S����{8�W�E�';!�I��#��T۶���;f��RI�#e��'o�또4����ZI�nm���6�?V��Q��|H�}������/����Q:�=���h*2� M�B�����������`M:ջ\8���L���G���׎N���[���W#����YU{��Ţ66����Z�W����<�/��j���2��f_�f}��T ��C��Q,�7��S]�y���c��1m�^q��H�E)���'���l(E�U�z�M�Q��5���MG'��g���xD�U�c4��3�q��?�ې�`��묽���p�4��G����w.����#��('v��2��}c���z�?4����}�l���q�b���t3�C���S�#�_O�}ǻ�u���P8����֫��Ho5f�I��q���ר�k��V�ƞ��y`$��,Vp�U��
N9 %�`	T3����4�?+�9o�E�tR�d�O^���S�w,F�u'p��{����ٷ}����m�-� ����~Q���N0xjfΖ�$��1p0�+��crZ�ȃP����-v-vIK-wQO[��*���LήLr#_���m��#�5�C��m���$�I}T��BԩI�����<H�[�;+[�0�L���,�ژm���OV�0^T�A�
�":�r���m�n`8ΎD��w.�5�W�L�#��·�V��b����p�q15v[�]��3����t���|��{�ڲ�O����˰9��)�n7b�B�X��E��(��j���=7��{J����]=t)�_k���[��d�s�	ۀ,i�;3!���C%��ˑOfR�8_GνzemVT|6�	Ѵ#���֤8>J�U�w�����.S�������+M�[ �Ц���0����;�Em���t8�M��R͙q��g.�n��Ǘ��,�5T��z�j�e�/t}�����]��K�
k_�����?�j|U��#-���>�y�q���m$z�����ϸ�b���j�f�B�#���b�]Z�6��`�y��}߯C��?T�4���:�Q���Y�4�I�7�&i5�=T9L����'��:d����
#�Ѵ�k��0�	�g}�G{7�V��8�l��}��~n]���v-_��cM�%�Ks~g=������P��}xn�$��o�Ur'���m�<k��>��ߚ��ف8�#��ר���[d@���9���ِ�B�Ӱ~�e[6���� :��:kܕ%���S���i=�.MX�n��\H2��Nү��ޓ%�Z�(��YJj�	>�ܻ��h��W�&N��Ǘ��>'������{��8��淬pFT�����`��~G�����6��!r�����s�5���Q�?��I��ɀ�hP�։t�&wk8#�4�Wݕn�.�;�K���Gfh�甓�e1��<�9A�p�w�\��/��r"�D;�67MC�k	����!���(TGt�����=���P�O�!C��.�����b%��N�al���,?�Wc-@���`F�'=��t�u&��Ѯ��\�#Kq�/��}�-�Gld��jjsf��	@#`d�Dz&�<��0k��\D�~X�5��䳚�^�V�1JJ��oE�TZ��\�0d��,����)���TM�A�KșR��݈7��Һ�@~z�������%蘾�0���S��d�>"���F��r�kU9un"�Q33��=_qe�v����!"�� ��M�*���_���ح#��4ũ.�s�ٻ��)�9�%�|x��>5�z��1t^ڪ����ɤ��uzlPA������n:b�$�V�0����%1�z�7V�<o��,4�b� q�I,8���f��d#Z��F�De�t�c���e3N)���������wnƚ���v�Ĵ�.�
XZ�����;�gM8�����-���+�e.}W8O&^\`��mѴsz�T�㒵a�b�禹մO�-u:kP7�֘��Uz�Bc�ᥔ��� W�] Xː�����F��|��?��:Wz[oBe]AD-�7{�/��^�7N�_Q_���he%
���7;D��K����+���uh*�)1\��-^������s���s�ߺ��Lv5�4 ����Z;6EWp�ǫ�P����F?�B��n�gq�N2pi��ibT��h�_�딪d�8����m�E��{'��8R	ƨ�%ߥ>�`b���$�-�p��������R0Ǵ�&[���i��Z��F�_*��%,����5��u��,F��ߧ,IQy�鿯�Z� ��n���d�PJ"\�I.�`C��R*��4Y'��5r��|�S�x;m�6���j�f��1F��;�<�UT?�,���j�/�@t�ƗH�HH�Hڮڃ�חү���3|>X�i�l R��ױH���d`y4�1U�@AV����4$(�N0�g����M��.�� 1!K�|O"Ź��\x/��%aI+D�
�)n����d?c))�5D�y�p����'�X؍J��E��\�?O��n�x4[�a�X�r	jV��z���>W�:���ܴ.P��`{K�iȉ����jG�c|�Pm���EK��n���M~nށq�������平L~�z'I9Dy2Ѳ�h�iS���^qѤi�����<�8����Msh�vI�{D ����.ڴ������I�Z{B�HR�οP>��$��jm	��#�	\�AH�&�z~?��A�B�U'��#M�����]V?�C�ECP��W�洍K��N�/�+	�u����6����0��0��g>��g���\��/��垚\#[p>�4�^��"������/ԡ,�E�s@�ϛ������ c�N��<��� V�tF,�ĈG�N��p�_�Tr�~�X��W3ָ�b�z�*�D�D��ާ{L��7�+j�s@r�#��G0傽=�W[&j!�&�A�k� ��Oeך�W��¯f���q݋/�ju׬B9��8�PĞe3E�<�y�sK��f��j�S��,B���
�� ��ˤi,��vɌ��iB���o�0�ٰ�ڈ����b�}���_J(bQ��j�f������Y?�3d�d�S@�)�}*e� �k��~>��72/~|������$�u�r'���"�+Jl����*Ŝg$�f875pjB7��M���zG�N�0*-ý �7�nU�u��FO�݄tҐEK}+��fXrrHp�؁���R�0�5�uh]�`��eD�[��PF�~�p�������>a_uE�p<�.��K?Щ�&���h
��\3t۱W�Ky�O#��r\y�lO���UQ9����o�r�����;� A�(����1�F���'��S�+��tJܣ��w?#:���"c+�mlg:�}�+�_���77�EX.*6T8����aVz0�b�,�e�~�B��	Ϙ���W�/������]�_LhmN��뜢���&�k�����l���FL��5���ۆn��#�J�i1oT�U�e��k���6<LWE`!PB7��d͆]V�y��d��	$��a��Du�8�t��������M7���{�e	=Co/e�����Na:J��x]���A� y�y��ds�|�)�����&O��׷������e�p+zn�S\�h��hP�����a
�ݺ���s�?5o̰tv���(�-y�)^����f�(Ra8bc��dvE��"��ڦ+����06jD�*��o<�~��*�h�fE��B�@�T��`���5!��Ϧ����/Ԩ�bW	�_�1���R��://Kt��LrH�NV��	�7G5�x>���9 ��]��xBҴy�5u)ȴ�K��;p�R��Vh�w��r���ɾ�_;U���*�M�ID
Qmxm�&7�|k�э{�;U�ԫ����w5��Z�Oso7�N�=��Z����5U=�$�0��q=���[~s4D�x~f�R�);�_��[���1��ڒ`=d�R�D=�zw�̦06��.����S��i�}�6x`���B�a��(<Gkb�f�Su�ɀ�>[8��b
��LAݗ�����E]��$��n��x-�F�7�,�4���z����#'@�G�pj�c8�C�ry���M�M�}���pg�_��L�mq����.�/[�7l���4@p����؂��	igb���&����Y�c�F$��[������E�����#������霙�)uӋEE�#�!F�N&�z��}V��
N�ڞx}�ߢ;{�!x,A��	c�E���E�wuI~f3bV�bc;̊U$�&C@�F2@S�[Lh�&�ve��R �{	�r����7z7�?�W��>CO��פ���1yq���$XZ�=���l�ꤰu��Ɩ����%1��޷$��Y0�"��/�"����YF|�;�r����la?�_��Y���Ur�a{��\.�u��6���^���t[xq����c��e�R�&�3E;���l����Ԩn��,ޝ��~�/+���ۤ���,�=Ҹ��&�U��-v��i���}6�ըp�h�/,��H���0[��o�E3e=�hS4G��2�,ŨǛ�� ��r-�2��T9�0�B�'H?:Ծ ��eXйZ�+�1�9?��\w��Sː���epwܡA�6#SZ$��헪���לTu񢻿֩��(��g��i��^  9�p�8�Ȳ������/(H��q~�[��:��޶׵�v��� �l���m��1�)�ю���*���ȉ�!6�����5.o߬���-N�շ���L�)���4�6��@���Enq�ߡi�f`a�|+0~�8��ir諾[1�ɤ��f������)�:���m/Y�]�{�|Dk,�ɚ��9��ڟ��nM���:e~�����[����'�q?�}�q�)Gw���d:�bq'a�^��FY�#(z�\M�(J��u���ۋ�h�.A�V1��ɐh�8iBז����������J2�o�AǺ@��_u�*��a�A���-�K��Ņ~_������ۋ�C��qU
JmsoRh�ه�d ��?N`Ky�3�K�:Nn���$����
 �\[��(\t�����@~�	]�+o�Dr�b�ä́﫛�O2T���1�:^��i���TȔ��'�������_�v�>�����S8]Jq�=��nG�9qe�n�;yhXc�u0[?�,�?����Ͻ��a~���NC���hs_� @%�R�0�)'���`Q��<���AuUs똇T��ǖ���r"7�b�����&�77�3�D	2Y��� K�D�v�h��σh�f*2p-.򼆢L�옽 2���I�A��TD�0H ��3�����"x1d�4dc��w��L���	TP��죓��g�yi�r�R:��MrM����1`AMA�,�����V�֐���I�}����`�[~P6,���F���c�C��p�S/4�>�z��Q�7�����{�t��zc9�5��W�I�F�u���E�����Cf!{��։���?,x3ć���Zd�?ߥ��uQ?uݢ�9�`�4��UH�sSJ{}�����A�I�P�ys�(APc��kJ�4����v�u#�|��
�B�==U�aq�7_��
�y������+:X��Fv��w4^L���-h/�HU�l1h�[�K�K7�aȻ������k�����\�X^�7"��Ǫ�!VD_{	���:����Zf|J���Z�V1���gKx��MV�����մ����x폼E�K]Ȁ�<b�N�Z:��ź�����BA�����-���z�67�����`�����e<���J�EF�H�q��mt�pY�Y�ݘ4 ػqܢER�Fm&�!{z�!�)oOdC�`!�S�Na�RK��ӈ�2Qb|�� �rT.���X�����d�ض�eR�I@O]�@���$ݞ�:�Cn��.���Nk���m��Jl� w��-p궹k��- ��J�l��L,�wa��ҭu��ﳠ�n[�X%��#�=(��*�H�~Q[$�g�P�"��m2�eJ�z��o�Ex�T�Â��:�yH/G<��������hF|�Gĳ-���"Y���ϩ�.�Xv�[�i��t���wq���=�=�_���\�,����@�.�y�g�5o�"W.*�����s�R����7"��8c�(��f���pCڹ�\O�t,d;���t�n|P��R�+\�3kD(σ�x���쪷���Rs�l7,?�:��o	�Cy4%��k��B	�)ތ傣3Zn/ɍ���\~����|����	���<.{�<b�O+j,�3�� -������|��'�tٻ�K욫�u榷`�!� Ѯ�p�,�����8uzp)G5k����og��~�.��5�#4u^��4�Uǎ����e��h��\휷�w[�<o�80(�o�tEd{�W�x�\?oB-e�jdC����Ζ+$Vf�N�r����W�ݧ�*5�'O���n����,��� ��%Q��"jA�i�����r�`ϰ[�� 0 �yV���jpD�q�حa6�K�UD�������zg��p��x���睟�,9O�n��]9���Q����
�h�)$�u�_�9::�ū�)٘������*zS&����t;��Ӥ��m���BX ��範k����!�Fmr-q��<�?�M#&���B/9`���~����u���+[�0�f�l\���J��|~S\�\r���_���p9S�}H|��v~��KD�ۡG4U���{�����kg�+��Ss+l֎O�>*�CZ;��B������A��m�1)R�BI,B�%��׮��"��9��u�^1�M&�S
'OR(�Z���Z��v=ƈwE�����5��׊��D��п�N��3����Mu�M��lb�E��N����ן]/Et������`��"�|TF�N0	g����Q8���	�_����#�K��W������:_��I?�	�a%XwTV����
#姱
=��I#�sGm�"�~����V��d��Z�ş�6��
���;l�6������G�J�X~2�ۗJ�mz�4�|;w�s(�� �gC)���ANg^8�^<�%�%�k��6Xd��E���Vj�N�A��my�M�rk���������'��S�鲾�6=�D���ĭv����3�9㚽�Vu�?,�(�)�7ޢ���f�0�'�.*a|͝W��w��)�[I4�ȜB��j��ЕX��RT��� CG���\|;�0у��h��G�TzA�̒��Uj�^�eo�uD�q�t��4*���a��x�L�q� 70�k�'L�����L]��\�mZɵ�V�����V�h.��z�T�-Vwf%@�����\�X�x�Z�A���u�DQ����{i�t�	�~��ˊ5eYZ����ɏ�6�7�6'F��σy67�m�؟}uu���CR�4q�Q#}E�VO�K�4'-n3��n�.���[��#A=J�:�q%)��!*��q�M�b���Rd��}���#L���B�Z��V��5h	���d�����k�_%>��n������W��S���dF�X�{�^��M�}T�|<��cR C��qc��2�6_�clB}�:3�{݃)��$/��!&C�m��� _��C�G��k�T)�k��{L�%�y��4�7>��,���b�������� ���|��ϗ�sO���H��~��G��ͲJ_K�M��V[n���_�a�g�om�V]��q���Zke-����y�"}c������֙��"o� ��5�>צE?!���$����ϓt�ԩ��/ږ��z�-��L����ݜ$��H%����K)�]�Z��FQh(w	�4׏+��ݛi��~�#��^�*��+���2�<�7�Ym�g;Z3�!iC��tb����N*���Zeh0����J�@�Ǹ�ȭ�o�ۖ]l�"�S݆����u������M��w��	2���kBp�B���G�oo��{;oc8�<�� ֵ����2eD5<�S�0W6����]ao[���2G�/���GA��1V�wM���8̞ �8������`��IӪzT���_q�]��ڷ�T��Z�8� �Q��N3�{+7lHW�:��[ԫ��F#����y�g<ڻ��' GOb�g��R;{B���$�Hc�co24�M#�T���|�6M�*cf.i�1�ѪT'��hu�7U��s@_菤�d`IR�$5}�\v��)�˅Qv � ������"�I#�`�O;E�X�����
 �JP��x�1��d�Ĥ�`k�׉��̅R�'��ґ�U���k>Z����aE�9\l8�&2�t�*����)���/9�C?%��$�m�G�H��?R��{�Cq��B��D��P;;�/�
+v���J��������g��d�������wz��Wf0��;T��P,7�]��d�	�2ajb�W��D DsB��d^���y)���~=r����ٕd>b���� 53��gz��\�U���R��Z��Ha��w��N���$�Q�c5sm@:8�hGP;S%r}҇�g��|�*vf�'��m��ik5��k	�89�X��c<3#���V��=�^?���5�r����܊Ξ�x:p�r���.�+���m��`�t.�7��&%|���k�F�p���e
�r�����zDg�*w�*�M`Vԋ�Hw+O�e��3����d��
>��T�ͷ�֗+�e�Fv�]�`��맴XWU�����~�+�꭭�}�
�{M{��
���8=���"�R4�jo��1�׶~L]�3�U���C��fN�K�jՃ��W ��)W�Vn�v��--�E�/J��������s��{�=��u���5��(\W��9U�YR�����b�v��ܾ�f��0��\3uh�p�t�/�ؼ��h�o���	`�K����.�L.2ٸ���8fd����H~c+n�Ѽ�{�_%������}�l���ύގ���R�k���\|2VK jS��S�U�~i/�~W�I�?�+�%ķa�y6W2�}깃A_�Ǻ��
�A*7�y�4|k��A�B��EH)��#��	1&��_����i��(����5�kc�J1���Õ�Y�W�EȒ�?_[?L����b�����D��$0!���U��`�$1ſz}�cUPך怓mo��,*����j�1(�6�����R����G0'W7wO7�R��,;�'tPĤ)����k�
�1�v�Z�A}u�ń�PM��Oy:v�Sq�H�a�5_�Ӷ�/,	9��=;��k0j���ډ�7����B��*6<B[%듦YR���vӶ-�uĉ~��t�1�$�gkNa/~�	h��ձ����;\/���?<���S������51�n氨V7S��5��)�u�b��}�<��e�;�p��xq����-7������\���.<�S\������.�&�f ����3u��J�3�#� ��.�#6��u�Tt�Nq�Oy�A�Ϙ(^:>�����C{�'R��Pp"�;D��DL/[<��&���k���=[uq2 �%_�Z����C4�G[����'��B�@d��o,j���Z�?W�D�F���YS�v��1�801C:�<&�riӪ�)y�?Up�۵N$�)S��'�r�nR^?8�%�8x<L'zF����^<ܦ8�\�W(
5S��H-��XUl��j7��w��>����$z�l�Sf�Ae��|�s>�`�0�7��Q&!m�;kT3��{��Dz����%��������2��Q�:;P�M߰�9 =�b/���w���Z]����>I�Xr51B����¸K+�^�P��&�}�Mj[ԓx�x��G�˧Y��4]یx��4�����$���E=���덦��L�xX��ң�ݢ:�XYSj�*�O�CbX{Ǥ����5ϭK�3L7�����Hcb[�H��ʅק,R��`�=�N���ѐ@�6��w�}J;�XRE��huB/mX�m�s�������r��o��r6���2��H���V���w�?fgs�9�3J��^�r7)�v�|I>�vIR���8}���P�h.!�g���y������X����7u���wT����l���T��)H���c�Y�39Bأ���]5x�ʞ2?�Z}q�� �3�Z�j��H���2T��(o�1��F�M0j�G�*۱:J+t+���X�mE�d��;؜gܿyG٬��.���o��x@�|k(��?ǁ,�F.ی"6G�����0�Cg��?�z����b��*%�j��#��D�l��PP���Kᢟ�ߦ��E�KnVw������cVPn�B0:���Q8>�}�e�SV�P0�-HA_����J�����/�aG��qn(�!���%�ѓ4����!^y���|�ˀ�]�E�'�!��V!2�~KcS���tfc���%U�2u�c����t��'4uA�%��F��A��K״�az$��]ɫ �аv���3Vk��ix^��
��Y�	�zm����0�xi�UF�.S�=*kW:[�+a��ل|�`o�^*�'Mz渦�z�F�w��`�����{(BKԾ�L}�:z����c�~�Vw)�Y>���h�Ȕ��<���-�by��{^{.��5��	�K=�[�ީs��v��(*�`z�������]����'�ה�x���ru�Ơ�P��rx�.�k��XAc�(Ѵ�8��?���]�9Bz�,���[<�[<���,��S�V�Cv�l�47��`foI�Ȋ�3�a�J�0�:��n}f�#�/A���@0�Vj�y�6�S��T~9	zx4�[)uM�a�X�h-�.��d��#�P�ӗɗ�~&��9Zܬ��-B���;O����n�6���3<�*=&�'�'��xTGc}\��y�SŴl�3���ϟ���ēa�X��52 �D|T�H��j�v�?����;j���*��m�q$wǥ�u/�Eg��דvt�F�4�ꣴs�5�NU�3݉��6�>>���q浢���dB���t���=�+��_�p�#v����\|];&}�g��W�`�Z�����C�f֔m�XΜ�h	���K�`5	ՍS�]��:�rQQ�ym{cğ�DQaڶ�n#��(.�(p��_w���8WB�Y�.m?]�S���/j�w����?�O,�h ~"��s3%��j�� |j��.��L[n_�Õm�p�*i:�>�����hq�X}�Ѭ�`����H7���5�P��c>/]�$JW.xr
�]Q�K���H�&2��$ud�^ҊB�j�һGmګM4+�=&����V<�hs�?a�K{�9L '~=�7��d�<�i��ܫ��$z���*�I�%1��,&���R�z'���l̨�	�پ�0���n�t���_� b��a�{H�!������<�H��u�m7�vu��Y�c�l�m5\�����;�����h��?���ȣ�m��L�cDV��䷯oS�U����m����l�e�2���k��[���z������ȶS�n����4�Y�Z�0{0�8L����1{Pƃ�{}'��\G{:�ʏh�_E�7Y_.��������DIx2��3-��#K�3�֒�د�i�w���Qdag.F�'j��Nh(r	���{8fY?�v����>�?��9����^N���͢"Z�;�.���|�g��?��F����hft;���$����哶���`�e,�ȇ�)�/,*��ɞ&��dX��"Y�Cn+X�O��$4��x��^��V���&�ߟ��� F�?W�F����S&�������<��h8�ǹ	"$��P�6�Hǽ�Czyjt8����>K{������p)o�9a����U%:���L�;}�-�s���τ��ە���	ф��|�:bZ�,�l���Q;��4D�_�绐r��Ao�3G���:|d���M�M��@���|O=>&N%�ŏ�2���k��Aӽg��[����SG�<e��m��!��M��
"T���+��T�N�F�U)���/���@ߙ���+�"��
9��c��^�|S1\J��f���j��-�N�k�[�C�����7�e�|~�Ͻ��"���N5�7O�#�� c�|Mq�51����	T�k��g��ӡ[G��[�H��#+f��ף���AM>_¾�����٩��jxZ�;�?z�ŶH ���.f"[i�٦�
ӲxTIAG���k�X\�K�-���J{�����n�:��O�:0�k
�'�Z����a<�ĕ_�	Q-ͻRN��Wq���V�r|�PT6����o����7�oX��
�d��`ձc��	Nvh��gq@�q�,�O=<ASwYo9�܉�8'��Z��-,1�?�mk� � �������wT��\ַ���@�FgP����ձ��bk�6���o9�&R�8k1&͋����>c,������0l�R��=��Or���	P\��G2W,��n�y�G|�:P��`2�ūO��"\&���`6��T�CI����z��O&��R��A��Bİ��(K0�_��wT�_�-� J������;(��" D���K (қ�t����{o�HG"��;	%H�����;����c��c$��Z{�5��s���>��Mܓ�|�F�ǹ���OH(���%,����|�������7a6����l���`��"��p���4�0�MjW��V'�f������̉B[_B��Lz�s��R�s�a�	�k�צ���V&�̰�к���� sd{
�{�+��-�{��^����W�j>'�E
ڠI���_B�zl��[V�!�\�:�[�,�����M 2`o~vL���~2c�u����`�������0�%��ν ��Jg <���f�h:��_��)�.ZcozL�Zԥ���me��W�S�l�}o���k�#�_��vy��n8�2�^���<�Ŭ�<��Ӗ5H�<�>2�-UH���� �O��pU\j�P�Ļd�^���+f:�剺�և]�$��~�b8�������S�I{3b���]B!a��tÉ�88O��ǐ�B���qc3��q�Nŗ@���Iҭ\����@|���3�\B���-w;1�I�M�۱S۾��sU�����Anȷo���ά��.�O�xs����1�#��jo��$�~��.{㌘$�ML���`��V�Ȳg*:S�pu�5�eE�W�'w��K~�U�S��P2��}ޝ���9�~ƆU�P�D��%r�,5�B��ݶI����>�&)�N�9�E^7:	e^!���#̹1'��lv����>B�k��t,D��(�D�$�:2����?�t�w�,-�`]��7.�=9��k�"�� 5I[~h�p�^��8�]ӝ@9P0�v��� ^k��i��Z��E����Ý��2�&L-r����ڊ����*V�$z�#����z�dNuc�1�{���!������(n?�~x�יٟiz��W.Å�n1��M뾗�K���)ݻ��`C�.p��q%f'�m<�H��/�e�E`�Qe�l?'����.i�����C퉜���3���tӁ�(��2�2�oiˎ�I��v�g��\�����F�T��0��S��/x��d߮����[=4=�(ZBz�e�w�BF��y�4i�$���<m�����iv2�Ð["ٝ�"/�	�C���K#v+Q�Ń&��
���/s^�z��;���6�d~�ī�l<���]����V	`��%����y)>H�a|<�{Ûo���yR���H	db�� e�w�O�Z��$���P�"یq��.P��ܲV�JgEh����z�U'�Վ�Y�J%1I'<�*"�e�/�M(!�{?��?}&���ԛ��Xu�S���8G����+�����YX�S�L�f5	���`}���a�]��3����Y�>6�0�0y��:t%˾���ǁnW���Â�<w���1�oT<#��_/	��-v^4��q$�	��Jsm�֤$6��;���K/sB��p{Kò�3wVՍƤ���Hu��=��۷�_���_����j��~�Z�x\ N��E��E�O�ɀ��3�9�d���"_.���jH��/ߓ3K��貯|2�� �='6Ĭ�C̿������0����tkh~��ֶ��̧�v�lA^���BS���R��q��V�ust�/c�py�('/�so�9iz��5���C�s�x�%��MBP�"��t����Bh]f�ξ���PkI�P�7�C�ۇK���y��~����W���f�n�c�#=�td�D�fi~�x)_CTv]�i҇Q��:/��ƅį]�~��?z�1�\�~�Ɵ*<c�]mğvM/����ÿo�K����F�p�"���REo~m���Һ���>�b�����o^y~�胢[	ͰM�	�^�يS� *�P����IĄ4K���ÅR1�5�!Z/���4�{'��}6�)w~l��|�s���=��!���5?�b�.�J���k�f8�_\�n�L�x_�P�������9�D��+m;�]b���ND5abˏ`�;�P�|}}W���3Z���D�n�~y�j���K􊏀�K����)E9�ˀ��vt��lC,<B>��9DA@���Z}���o�/�$��Q�QU���~�%�5�t��ǖ�ͤ3��Em���y
��[��ϾH6#Gz�Z���Jz�K��?�b���O�UZ��\���^ O�A7�Wm������ԺCm}��oHYi����@�����Ϝb�����T����U��Af���>>w�����P�c2Z|�Y�C�r��dZ\o��Hnx1��a�=H%�|Cz�̹��E�(�r(c�5�vB"�y�X}�HMy��t!�|ҷ{\�n���yYk~}��R�������|���ܿh�������Q���t˰��;pCT��u��GA�7eΐ��נ>?�Oё�A��w�Kf���������,�O�k��0]r��%gр���}F�\�Ԧ���'��ٖ�]n�B�g2���r]�ޔ˿���e���N�2��]t'V�ϼ�j�I�qru���ص��m�Za��u��������^'�����B|`���ȳ=�~����\u^��uNm�W1κ�>�&C�צ����8���?ܼ�>5��4کDw��Q��__ ����6S��@�V��#@�G%��5q�3�K�M��pyG,��t����w�\;��;X�=���u��
I����s?[^#_i�9D|Cð5�����sⰪN�h.̑+�S�㛹:�	m��|<g�h-#�����Z��G�I��-j�Iu|�Da��)V���a4}�U@�V7�TńPb�*�}���p���h�n���}ERZ�N�B/_��XK8!�8���K_�pi�������ۜ7у5�n�eڦ�h�`6�լ���{7 �u�3)�f̛�1y�㭖���5tS��98�N��2���6��^�w ;��*z�+0[�U����2U
c��v�&�D��?؛�oљ��R����A�	�+8�(��ޢ�Qh^�R��Ն��y�U�L�}�z��=X��9�Ke�R���b�����<y1����1���^�n��2��F�/��rJw�|\��>{�v+�u?� L��x�5���_��G�@g����.h�d����]�A���.%���L�a���`���q��b�pf�v����2�����SW5: �g�x<�ɖn,�Ѝ�[�d͜��a!uo]�s���f��2R�Z����z�N�p����8���V����+Ɇ9&�d�<,w��1CǗ=Gn��=Z��x�k줽��}Jg�aUF��o'��*���~�3��2�^��}r��%��'��7�j��?�ZZ�'�������D����V޹?�T���$�sX��~�� ��=g~��ǽ!�.^��]�aO��|��@�o��ٜul��A�"�|��%:]��)��3�u�ƫ��y�VN|Zd����<F����~��aT�M\��K��;��NG��(�ߞ�hW�zFS,ׯ��_�2\�I̋�ݪ�㦯����fZįk\�!���M96{7�Z��H�W���N45	�:Tț�/Ż��y�1�[���E�:��9����I#?�7*(/9���<x �/�gj����]�����8��h���ҤԮ��b0���S�~���?u����m�MXG)��KЄ?!D�.a�ʗ>OZ�q�����Qh)>��8ִ��veѤ��څ�\�~��������[���iL����⁫�
������uu�;�&��h�/X��6���P���3l��#�����G�
�iT��(�a�*��Ο�b��aW��5Uy��R�5��2��!����.��A��ù��&Οx:Ӷ!]I��#���ǰ);�j�&*l�}8ù�U��b��-��~������?5�� �K<g�yDw�غM�@��u.׆��-9U��+%?~�N�o>��a�C�?�O8���Pa8.�(�^ֵՠ#�ss{?��:7�!w	>0�)j���T��gi��fgP���pzu��!���������A �����S#�}ᩴ�pJh·���/9T0�(>!QB�=.\��c���4�n��Y�9x:�L�A���(3],$.��u��x� �W��0���Q�}\�����{;guq���zB6����v�#e~��h�~ћ@��%@v�\ü�q}�V����zk�Xޟ݀�����g5�����2�-ܩߧ�*LB�~��nB�2(��>yU|O��Y}����:���n�	�T���U� FoI���8q��{ۯ�O)c�|���i�����tY9�OG^���;��N��E�5� :\��?B⻏�w�D���<���>tSCS���e����qU�F�P�����iZ���p�XZ��2����֣F�u��6�Zg5j��%�Sf	����@E"�_5���h2�/�\ (tAؾ�)ŋRk'��﷜�1B��}+'� Zy��Uҍ�;o�W3>�>�$8!�(l�J	�xx�n�N.|��ar{�EF][���\~Ž�x?r���#�)osd3%m���X� D m��3�qЧ�`,����ß����N�A��r��lR�6�r�-��YƔR{���h����_aQ¥�_#��4I-6�����_KV9O��v���+��~���`R����DO��N�|#�WU�+��4����x�RN�ɡd����A��6�̽\4�K��5��D}����M��m��|�i�R�8� O[��ͼ�i۔xps�G���S ��̫Xv��	}C�?���}�O�J+�P	%�Fn�ɺ/���*�%X�\iݰkEK�bp��������F��^���4^(��;Oqi��Vj�Hgl��7 �ʙ[��/r�]���
zS�ss�=gNu�T-�e���k-�#�6&|��ݚI�љӃ'����@n�Dq��t"�,T��D�?7��コ�����kY�gM;�V�ΚW�pݑ���,���+f�	�����%��86,���G����	V������JM6���gѺQ�!D�qyT�s6����������8�O���>��Dɐ��髳R�4Yi<�1c�iI��K�O��g�z5�z�x�����=.ݰS��u�l&T������zH�6k�8����U�����t�����1	L����W�o��[��h⒥�8d0�:jl�7B����G�Oy=y��/MC)v΍�n� hK[�p�������%g̎�_~�G�vu��=+n {�+ȇZ���ީ��rQ��<��u�A��7<�ve��kw��f�\�C	1UsTz��e;V�hz�1^�������Z��Z����Y�it�쒏���1�ޅ�"]����U*CV����#�E]��RR��j��Ǖ�j�&ʹXj�"#[�����&WSU��pH�tԼ!F����'dV�)e�\�/�yuѐ�d0C�2ip]�g�ߚ=�ϧ��$|�ԑ�Z�\�u�/��+A�j��	��~�/&��k���"��bOaYpB%bF�s�
z�Y(d3�~#8���+��� ��1E�� �[�g��&����ȁ�e�� ��xrг]���svYT��s��X�V�͵FL��N�Vd$~�M�~C���s�.����iKD<o�@�˨,�?ֿ݃��մv����BM,Ks�Ve�c�%O�7d�z�>�մ��9/VcClI0�p����j��ǉ��2w������q���/�M�����K�Oy,����r�&�c�k#�l&A]�:}+�������:P�+o�3d�:*$ۥ�nU�!���f\�ߙ���+���2�����UM:w�&[����텞KY݈�L'�OI��� z�U-�lS��&�{���!�u�Dd�2:��Ĳp��y����+,W���+��R�.NQ\���î�	�Gx�qun�T��g]�(K9�X�9�UU�
�ä�� v�G�7[O�H�ހཫ{=�73�H�>�gMO�Mp��� j9e��tz�p�-!Zi!���Y�O��t�u�9o�����ݹ�N���l�:sD
�4��w�~W
��AVɯ�D�� ֻ-�L��GOT��se��fȝ���l��Tg�PI��B��k&ڎ���W��v���5�qz\�u��C���G��	'C��2{7c0�t�lB�{�m��
-�
�Uw�8e΄�{�2쭄��n�XWFzK���] e��$�o0?{(�`f��8ȗZ?Z7$u6���o:��K6@s+�yx,V<�|�b_���	�:�(N���\�Q3�Ӕ���+Y��p����O�d}����a6�x�"A�^����DW5�+�9 .�q�������!Ѭe��ʇ��^7�{��_���@����E[H��Ĕ<a��
��$�_(�u��B�Xݏ�J���s}cq�i�J����~�ׁ�I ������B�)U��<��8j�d��x�$��|ױ���+����건}k[���q9�>�9|��3�4k�C{ؑ��:�����V�<z8A�[�VS���b5�ٺ��di��~�U�B��	>��dGМ�~��-y+��9�%W���j�2]E�}I���>�0��W�-�P᱓Ice,�}��r���*��pLV���\fX�#K���	� n.덷SW�$g+@ S;���=3�A?��;���p^c���|{���i\$j2��F���21z2�͹ ��ye�g�;��� i���*4���z
���m�&Iy��u�'�p|�^H��L:��M��ļ\n+��t�b�w}c��|7�,Ѧ���G�Ƶgј�)
y��dM
��f;W���&��:N�rv��UUΊ~ڑ�~��:����	R��mY�#rX���(���)�y��
��y ݧ
��H��H����)�����␩3&"*fM�Q�f�80�]�ˌ���8��/�Ɇ(4!���Q^!���U,{��d�ܚ��N~�D��f�nX@��c3�lYW<'���嬛M?�S���|��gl�~]�a9Ƕ�ˤ2�Ʌ�d$ۥT7W�L�>�--k'j�͚�+y���(z��z�.~{�N[ho�Ā��_@P3`Z��qC-�=�\z����G�k�l1,\W(G/A�����d�H�K����R;���-���i������	i���#"�v��'���o��cJ�kH�L-oC�>o���j/�%2�t���Ok�����w��jK1C�|��ɣ���/���C�OL=W�nX]j+�x5��>�Eߙ�Ϲe
����N�{��f�)�,� ��rh�6~L�FW�V�a�oZ�%�Dշ9���	��uY4Ix����� �� 6>Tn�t�����E�!�qE�V�6�'��9>خ�w����S�����ǵ��P�8��A8�ʘx���-+4�y�.��j����Hd?��C�y�E�ʉThl�BP�;� ^c�J�c�Y���WHz�X��p�ឰ!��#a���g�Q�2�n'w~�~'v���w �x8�h\���X�ڋG��-�[W�i���H��g�?_kQ#�`b�������?�%5'd�@����sH�9�4�|g�k:(K�hbPRQ����s�A�;��B�;p�p�u!Z�~�=�a����DD�v�	�_'����ܞ�"��r�F��!7���h�O�ř�o\�d�� 4��s{7C3�� �wPu��93��xkZ1�#�.ѷ��Y�J\�ɒa'ϯk�d-�8���;�zm����Zd�f&���(3�IЈ.�6:��X� ��� ��_��<f>ɉ�K)��>�u�i]��s=9�l?7J��y.���_R�����9s
�获s��^�p t��PY���N�*�?T�� ��{16hG�x=�"�_z����>�X0�?t��
Y���[����O�d�:V���q������Gb��5w'(PYFb��Hw�u�-]�Fg/N��!�� e2�΄������,U���(���5w�Y`Ah�M������^��rm���CV�	RjLqс
qoG)���֊��I^9)Z�_���D�p�����ߢգ�9��"�J�d��9�GWF��,��=��5T����'�Y��1�3,+�l�o4���ϏHZ<��p�Ⱦ5��ӄs�B�,���^�!���+�r���^t�� ��;ZD�2�0�%��쌻�=������a��@7 "	�V� ���v������9����Q�q�S1o�]|���nm��䭌n��'��g�=~�x[�8	"?�>[�@�t�C�س��Y�\����E��4�Ǜ�V�T�С��T!q�44Ug���d�� �P��P�*�W�ـ��,w�A�D�1qC-���pc�ۖ�?ڶ��=�,p�9���;�
�E�;M�t8/]bo�x��_�ѕ=B���?-�Xf��[�І"h����}�>[�SSvdt��D��eũ�V-L��$��@g��l@���!�k�ɵ�	 ��B*7��7�,#����N�/�:�rk<���ak���$Y������`=MK���Z�"�o�";^	U�ԁ�
|7z��)�=�f��6�Ű���sQ4�en�I5�o��X
�w��U��~B�N�U��X�s��\$��[ߌ>hR��,�c��M�G:Z#��׻�q��W9��&9�
R���~��z-�;U������է��������z������I�
]V<�{�k�8�kϩ:�=�=J)�\�,0�Dq��!01�T���̞��2��(	���Iȥ�*���vBWѷ�RIi$�����>��h�h��×�������W�x��,鍙g�$nAC�4&��͕��{7�ks��E��\��dJ��M�x�����_c�����J���޺�Q ��%������ء3g؈����ŗ�#�c���9A�Ն������,��.	�^.G5	�]_��&��i꒴m�D��.�D~�r'���@��Ϙ>B-��KJ�*L��78���k�-Y.�-���:�KFfp�a%�ڈѭ����M)����7]���3,�|?����|�!0��-h�Է^F���a�=]�1�ί����FJY���~������d�9ʩ��Gգ��X7^}��CK}��sm���{����^�j{����;�����&��[���l��{4:���]�hYcm��F��#��vp�f�pcy	|Jk��i�;��A��0�� �,��$J�a�RA�ޗ���V�'�Ń�n��T���j��:X�8q�,f��Yܡ�����G�D�h���e�e����^��ķ�6�3e����d0TT�P�6"�.�($�U{m&�{���IƼ���Zc19�i�����z�p�T�'4ٳK����f����)��d��H�b�,��=��T#�)�^�D���1�91	���c���8Os[���0�'�b�nU�_^'O�m�uI��3�0 ?�*�
�C�n[Q|V[dv[�����M���^��� /��f(bj�P���ŧ�t�����}�!�S�^��oϠA����6Y��g_�8(k�nL ^��T�/�3<���)�<!�2�x�.���6OH��u��v
p9o�Pq�-6�ƒ�\h�1���q�����9�]�D�I�^���S��h�y97�A��ѹ*�R#����i��۸St�Hм,�j����YS�ժ�51�](@u%4��N�G�4�O�^�N�LB��3�e�X�3�ħ>�5����x�Hυ6`tPJ�%0-x!�)���ӻMf��^-�bM���Gѧp]�%j(���?��ZLI��N�ڰ��{s�h`�L�F���~e�h{����S�d8����:��.qEteޒ�)��Y�k�&ج���=,���M���>|t�Q��GK��uT�[\2V��D�!���%�J�~�F�<q�d[7��F&<~��S�4���FO�%��x���3I��ކ9��;�t����L�7�d�v�j��rl^�qn��Y�*��D�&�1��^��}V9X��K��	�9����v��߬��B�����N�^���ua�s�$��:�,p=pNf�tZ��ƣ��3�;���6�	�Y�eX[�i� aT�~��>�#z(���-�De�do�q,;˵ܷ�Wd�.�&��t�������i5�G�M��M�b�%����V7���\N?*s�&R�<���Ǫ3���Tʃ�/�+����f�Q�&
d�>7����C�f=%0�<:���7jiUz�=Zby�X��(EM=쿵��%�[h9M%��>���<��B���JF��/a�)H^�2NfX�����[�_���r y\���e�Y�W5�Pi��z͋t_��x^��J�!��i/	�����j��C�G/��9D��8��{�� �4R��.�������u"��.媍Ѭ�����R����aC
¦�5��ښ��qkt����N�����s��7��R�+	s6}�pt��H+"�x�wh�ӗ)\\:`��cX,��ꌸ�q���Ͼ���h��O�.@Ȟ��
Ll���j�;=}��c�>޻�P�;"�x��{�v�؝���v���u���e�5jS�ߒr�6N�4��X�@���>�������My���{/�,�G����BT�ͼ��\ju݆2Ѫ���"�K�Xd�o}��#3�
�=k�#O~׌����-ʁ��07��^�_ �uU�j��):ߩZ�L��������^����ը�ϼʰ�D/�_jp}b�~	���ıC_�=Hy#oē/�������lk�#}.�!�?^�F8�v�pd_ Y��#���oO��Ii7p�M:�����/a���1�(���A�J���h�M:�?\ ��4�WRh1��q*�K����i%_�c �"E�]�������Yv��R��i�i}麽��Tl�b=����ӳ=��!V�������D��*�/_ ؜�dC�et�Q��x�NTW>+�����y��Ϝ]��s"ۢ0i�RG}�����R	^�`��,�e���K��+袹a+���C�ϛJf%�Κ�r�w���I�M�MD�T��!y[Xٴ�Y;�;�or�\gӋ]�Z�k� d�4A�9�o���ʻ���R�?2����к�����;�N�W�ni�C�i7�qq(7-�a��_�´��͂wՁ�,�o�b�X���|���k�X�T"=M���r/q�)c���'�Br�2�ղfO�NgO(MYB�d�_����Z��Dm��{^l}C)�H��ň�t������3� v���4cu|��wb��G&7�B�[r�dLy�FgG�ɩ*x�����=9�(���9U:P��.xT��%���7~�E�I� �;�rFf肥�Ȏ}v�3BK<㔋#��pg��+���$gN���p�N,�.�Kr�f_�L��i��&�e�92Z6e����	>z�	Ʊ1]�e�o���RO���Z`���6���[��cֳZ�利(�����r���"E1�[�k�<�U��%$�{�X�nl�K�gC��/��S��p#Z$B�9��2~��B q��nC��V��R{�5�I�"��6iP����Ɇ(^
�?u�o��p��՜�n^'�3�>��b�6=���e���/��
�����-�C(�m�ka�Kj�0��W����g�Ӷ���1���Y�B�ݢq�o��G�SmJF�Z�2���7jY>=��{�bC�+��ce���֘y.�:�u�X1N�esu�u��Ө�8�����-���ر���"���78ݮ����h��qj���3��	���q��^��[���z�lJ���>�]��S��zA�r��,ᇉ�r�������陓[?3��[#�7 C-�y�T�#�%$G��'Rba�=h���>y����fM"X���PUW��b0[�G����ɇ��Gr�R�E���C���u�S1ta��l'6T�s�0�gM��V#���䚮L�c4��~�O��U�#��	�����q�Έ^��d����X�r�`�,��^=����T�K��N�吽�r�3�@�R�^Ń�_�V����z�Ӯb��`t}�%�}�ٺ?�� ~Q�Z>�a [��ی�L��1�n�j\ii2o�`������_@@��.��+l����t�R���� �Q���<V,���5Oe�;����p�|&=�nX��'O8Ƙ�л�/��<��������hބ��,��C�H�!!�^�G��ۮ;��J��7��_7����g�wv�',VW�J�5�.�Y��wǹ�P�7����e'w\�����b�����i���b��s�l=���P��ZD&Z5&̗3I��>�;顱})O|��s}ǭf�[m��r��H�7��蓮V*y?�q�6����̇���5�d]��gq��F
��|k2�_C�Ɗ��[�pccC�!l�۹�zW
B  �4ֆ�ו�ol�47GG(~�(X �%�MM���Fv�^�c��g�1|ۓ�'+sr,�s>���;�-����h�������%~s)�w�Г�F���;ܗ�ǅ	9r�� ��
2�N�aň�E�;%ͥ���L���O����0p���B8����ꦉg̋�2�v#^��ԥ(0y$}5���˛�/�L��LzF]��1B�F�*Gw�UQ$�&a�_\ ��wkr�JK,-C� ��t��� ��� �]J�̤���*�hD�{�6:�:&_�U9���`����tJb	�N^&vf���)ٽS����VRl��w�����'DԹ����Ӯ��1.�dC��Z���K7��Vz�#|�ߢ:�`pW�ժ5���δ弍��3���G��j�� =�ew�����q��M�͐픡�6W;�L��]�_�c��3k>���;kټ�i��TGٞ���pWD+Q�.�	��UW"|Wn�x6�6s��I����%
���&���m����3�O~	h��=$7w1����9,��X�����^��t�eO���֓�!�]�7Kv�f�^N�>�#ᖬU���w5_��F��d�*�a�w�/R�uz�~�)>f��G�����@�*?���Ezux"��9D�,�H8�T�t�}�"K]
Ec���g��j�\voJ�&G}� ~;��M�z����[�ꕗ���$��n  Ǆ�F3,�I��w1��Mxn%1z�Th��0��'b�p�SO+�	�	.��%	�6�,�,/^zR�޳W��P�^",1V�ǹ�)�BMs[�;���/�������Z��W�
$F0]wU<(��4#|���� h�C=�_r�����6:�����(犿��w�<�
Ou�����8"�j�r��y1+�����j2�n�d�����"�6�I6W�7�P@�V�����hQ+�G�:u<��do�¨�����А؎)�ފ��� ����)Ô�@�YW�W��U���c��e"������p�8+���7�nx�51a�F������)N�Iz�hi���:�2>���ϗ�f�y�q?d<h����jk�7MlTm%����Z瞽y(em���J���sŏ����d�U⽻Ͷ�o���Qq�A�ǘ �T��~̾�pgӥ�}�	;K��s���ݜt��M��p���U���0�|O���U-�{��S���}I�+30���(;|Gu���Ѭ�m��2���c(G�x�"�P唭�&ѱi������=��OK�ƥa��Q@A5 =7�Cg.���д�8�R]���CαS�e�d���*���b�������t�W��)�Qwv���X��%o�4�f��:H��j{��h��ٔAO/�N�b�9�4�R"�����%P$kz�|Z���kmUՓ8�4G.zM~Rބ�b��៦ޝ�I����c<N�_�|��8��=]r/f~y#d�f9�6�M�e�o�s�����ʪV�W��䞦Q?L�y���tD=m+ҥp����[I�?���O�3����dd�;�5�[��"]�̞Lw,�+���.�Oa�%h*���`q������k���Y4�?Z�'�C��
�8��&$��m=e��S�9�2�R2������F�-�(��i��I�	�k E��r��@j��/U-��|�}��>�/��2T�-N�lH�Y�M5T�v<�lA�L�T�_-~�Ew�[�2l�+UӛO�4�����}v�^��н"uei6�:�o�W��/��d�����g/4�h:g�on'�j%&��#Y�_�L)�9�at��S���5�Id,��ɪ�]�i�ȗ�a�O���C/,mXkoK�8�H��,������G���G�$.=�ۺ+������P��t�A���,��.]{�(�8�CW(�z+��$ߝEn�%�'=�E��|m���&�c�~nb����Ӿ�"&���;�l���̐�x)4>��c�6�zi�(��is��7��*d�"��>���v��ױTN���	&�7�N"U�
O��:e������O-^䄽����5ƄD�.��] XVcF��q�z���M�12iζ\x)������l��֮V�n�8u�����@�[�zY�d�"��5U�-�āqqȀ!+Wlv�t؃���0�e�n/��.i!�Y$���DT�/ s�@M���Y���>:��͚,�`ۜ�_�8�Uw�ZR7iW��xS(A������j�$h��f��j�#��[7b�n� Z�<�ޥ&�54����=���٠ǜRg M���V��}V�z�m�] -�3�
9�;�p�/�0��hJgUw	�`�يp��V�����^KsfG�M��	��I���Nڙ��-���1�Z�*�h>\bL�����r��B۱��%�]���~������X�﬽z����˛�td1��	\ ��0� )���nsf��\0͍y�C�5w��9����"�<qq�K��;�]T��F���~�-��;��q��NKz˿񔤊$��^J̊��E�^�z4^�#�.\����G�R���g-[�o>n�jD�E�] |	�bw*�@_�+��PƧ�v��3�Î�!���ggy�H7�_5�Ծ��&d�m2q7e�������o�^ƴ�ٴq]�NM���[��CXEf�Ε7�Σ��KS�1P���� �K��>�G������s=<�u�WKD
GS�	���e �`܈�{�ɹؠ��P�������VU�e������o1�9�=K��4hc��ȯ�}�)Ե��8|�W�#� �� ��y��g�L<[]����������h�<�`c�Y''��W�A�������kI�#�S�w��JabN�/�'�-�8%Hddn��Ƴ�����x˫q��s=�� �??ML�(�r^UU���佹���]�#��Ep�LD�f��11N�:k��Y��I�2H`��a2��a_x�����8g�m�����1����;�6��L��bqF��V�Fg}�l�3�=/�oΥ��"m��*Z)ƞÿ��e�s`��#�KǠq���I��<�a��W��i[���k�r�0�רdF��wő�����a����.q��?�K��d�C��'��F�< pxԬ���`�g��Ju�;۸�ws  �-�&�@�`�${���]u�����6���Pq=J��Z�`�x���i(�ñ��/�j�ˉ�+�&Hi6M>���}�׳W�\�H���pnqpt�g{<�������prϚ[u+��`NMұ.�]�����gly�4��6��J��t-��?;��>|zbH����"��q$_sC�����1I�=���4���4�ϿLjE��9�z�ٖ�Œ��p=�w�+��'��]�f0D��A�W��H�ּ����F73�Ӂ7K�	=�׹0|yǑ�,�c�_����r&���=�:2�9�Y���|�������ԛJΕ �i��Xo���)��i�٘���7�bDo���]R^�z)��H��	747�$�!�F�d��u�T��hq[^W5M�,��Z���1�/�Q�����O�#]�rT&b@�.[�� 13o���x����K�����8�#��s�H��c����`�����y׋ٙ���so���a4�ʜ/�q���S���]7�z>G���\�w.�,$~�z��`iz�n�U���$�E_Iҏ��R�'O����a*v�̭�^Ob��фgA�S�̛�1_�,}�S#�Oc���'̩��A;�2��,,�Sm���U�Ӻ2��@A�u�����iu4��9���"����A�g��?�{�=�Q�C4��ح��'9����I�N�--h�'2��/Ƙ��I���K�:���춛��R��Rzs8�>�;!���H	��L��3�Ex�;O-����뷟�X�:�@�P��n=ӹiQ�-6=��S+s�=r_ c&��<����t�� �:ï��/���:��ʫ���d����\��������B���]�+���|U.�,~�
9~Ve��x�G�Hɣ[�VC��T���|;"a�$��t���Q*MZ��x��#O��U��+`��m�EK}�����y���7����PB7Q�2����������~mk�[ZJ�ew�Cbi
N���p����Iv��{vxj݄�~�?��搿۴m�YiCuz�uӋ2pၿ�qM��U���˽�5���Sw�'[~��us�Ub<���ۦd[����<ʶ��R��Cd7�%�� ْ��f$["�&�<�ed}�,��Zcf�/Y�k�e�c�>։1�N������}�y^�߹�����r��}�3Lo+f!?i�>Y���7憈l��\j��8��|��A$6�%X�� ?]�A������ƍ��B;U��k{��W@w��y���~<�_W�`�-�@�Fa�����Z��j��(���i2ҝB�Y�S	���&�oJ����Ċ~Y���FN�y?�Ђ�Nj�zv)iA"��lV\}�e5L&��]�����Q9��[��_4us7�Ɂf��b��b����hg�fK�l�u�h^{�p0}��i��YoUb�R�K	R�����ʐ�_F���ݚ���ȩwi#�MUED���Y	�sbO�;����.&���������p"r��ٴb[������V�7[����TŖj�O7	������y_�R����z��6r
�*�s�bS���C(IDG^�j�����{�܀��_�%������@��/$& ��|�O6{�����UFoPa��}l��C�T��;#�e�l=�2��i�� ǄM��~���.[�M���Wg�Ѱ���H��\ޥ�(zM�	+	Q�i��?�R��Y��Ct'��VD�{ΖD�B�mlf&iJ��J���"%����0YRQ����W7�XZ�S��F/ r����\�󓴜� F�7�HFe�F�'��\���f��ۏ��ʲC�ru5/����'���4~}�gL;<0��}E���&���AL]*J#�W���(r����4�K��g��\ނ�SL@:<���Y(l�Ɯ����>$���y��\�	MW�:d����sYfb��4���!���y&0�û?��Y�}�Q:��9�jRi�(*�@�B����ԣ8��S�	��P��$P�Z8���t���gTR9���0aj���$$֗h�����A�Ũ�<W~;�����I�I'��ʢC'�	x#3mp�3z����3j]��*����<�u���GD�Ԭ�-��Js��zq�*�v�� ��������Qj�	b+�kM���0�$򐳟U%ˑ5���K�݅O�CB�Q��%�f
�6Ș�hW(p���#~jG2���2��;�wcШ����lmy$ŲB�Ĺ�����"�z����L��Y�(� Aػ�CW�:X�::p�/Rݗ�������5��KgÑ剴�$� �oGQ+WL;[��ʥP�B�3�d�Ջ9{-s[5����_Y�~I�c<iQw[o�4Ey��!nv\�g���`g���S�""&�_Kx��ϓ�ο�L5��������u���DajM��#����S��s��a�[j(�Cݳ���j�F�L��9������x/ט�vB�@Ǽg�q�����!�c�U����*5���������2�=�B���^1���o��=.V��e���.ڙ�/�&�i~�a��v����rPd�	�0�1���q��.��n�\��m�p����ş�s}^�2$Y�N��6����F�/�ה����y�kv��	,��;�f"�6:����IȾ%hr�����53+uz�c�Z�2����#kj^��}�x�`E[�z�ʹE�.D��H���1{Q&�x��;X}���v�~.��K*���!��s�`��,F�X�h�J�j��V�/���(Q4��3�+xM��4~���n�ɂ�%:��PR�[�Ow/V�'�>N�"8��rp���%Rq�ZB�5���E��+�o���"qi
�ŭ�؝��g-÷)$�W�;Q�����c�2�2��|ǁ��^:�#��dc��8$���8�"�@`M)�.����I�o��!������m�=��E�`���'Y�����3Ȑ����
���ڍ�{B��ߟEP_h��>�n�8&�����={Ra�=Ժ,f{=$�	��T�|���J�|z
�_�pIL୨]Ύ��6�q{D�*�IQZ]�<k��Ag�j&�}$ŀ*�����?���F�&'Tscx�n[X�2D���l���0�`�o�_���;Y�;h���.0yS�%ػKE!1��������F��t�`hߟ��/�I�������'�E��m	���Y���Y�}�V=���bt9�i�S �\R1���|V������n���`���������f9d�;U�gmϾU�Żs%�-_�J�����9���]~���]EΌ���~ޮ�E����X-��?`,`�xỊ��6���&�wn�L��3�>KW�>��ژ7K/��)�W��?I�h�L�tx�*z8�;��'����;X�^���|��]n9X|�b�����5�%�"��dֺ��5���le���3i��K��Q�䦭�Q���Y����NH5�������s�r���F�Km5�rɽ�|�0{�F�~�%
vf,����f�:�U흗���#p�~'!ݥ���x��d��cp�����)a$��$��|�b5��v���@�r��-ٴnL>+V_�K OZ �\m�b�����zG����;L@l1�/)z\��*�_Z�f˂I䇣��+(9X�E2����Ou�~V�ur�>�c��I߀��Z� ���H�*��}�V|�ߥ��Z�H��c��Uq�9cX��os[y�՚[�IΎF���������~a�W�,q�Q��݌�&�/U�+�b�	�-�!z������/dE���D��VJ-��sZl���.���.��i��?�E��N�FG�T=�j�p�ތ�T;�F|�
��m��0�vr6��,-��GO.�x�9U�,����d������
?�P���"�U��A�`u�9~�	�%�!B��Y���!�3
���O"�6l�М��Lh��(�H�1� c���w#�Nt���a��>��)����RQ�A�pc�e]�Q��O�a������:-OΗ��kM� A���t���߱����ޔ��}���R(�pR�Q�[Jͤ�}����=!ԕT���?�MY���X����&��Ey������Le����]z�QF�^s&2�ͭ���{�6$І���e���F�ϑ�Ʌ㪳%q79��D��tݙ�Rq=�Zשs�w�ȝ2��E�(�f�~�o����b7�	�gw��Ep��8L5�P,�,3����]�?.}Q<z���W�9^�P ]�3ݭ�O�8LMmB{�~�!�]�L�ؕG��g�粯�d�;�0h-�%�5{��l��p��]Q������@c=�Cy��7��j)��yw!^��]u��'C�=�)�3�v�D��eyp�7�W<��h������+o�	n%�N��7��SrCg�y\��@��mO��'��f�?��3��R��Mܶ��#]���!��&��&pJx�d�KN�6`�����#ı� �K8��M#�p`x��N�Z0�Ӝ�\�<�!�U�8�u�@
�6}A�F���E\U��lr�A��I���K�5��w�UWn[]���6+0����'�޷n �u&H��G�&�4�X���"5Q�y������`��Z)0��LrO��_��Z)B���Яf3��Q6�L���k��/o��b�[x�|fa���i/���^�m�RU[�{��O={�.�
��f�����P�PI����܎�y������3R��� ~�f4�������~����u}n���*?��4�r�p̛@X��JÕC����{��T�#,8�B��+�P� O?�k��5q��}W�E�wL� L;=�U^�?б~yE�B��xk.|�-1nN5��q��Q��@��0�����~uh��w��\?ID���� ������ڤ��@073?'N&�>����*G��sߔm@��~Wq0m�_i+�1S1,b�ʾ�݁W-�3��Z�8�O��q��)��_���p������&�c\��}��SǯN/�[��/D?�J$$[�XF�t��o�7?!��i��^ۥ���c�������+ɪ/�.̼�$,W}%����}��oު���?��Ʊ�ǲ���'=�6��W�s�<:5�![/�틅�졹�M���wO��@ �w
b��*[���D�m ߋ;�d�;���P𰖴�s1d9��v������(5��w�ϪY�f|�ԑ��1��G�Y�3��PK   b^"U���3T  b�  /   images/b0310726-02d1-40a2-b36d-0772497b5f9f.jpg�	<�o�/���%)
a
Ed��IB�ƾk��$��R�0!�	ْ}��.�]d���fy���������s�缞s�3���ޟ��>ר/b?q8����
��� �@�pU��� n� �  8P4 )X� 6 ��:	�������D�������9��/�l �N� �A�m�`��rX�a9,���_Z��Y9�w;�e���tV�����������������������8KTXTTVXFVX���������8 P�$�=+a`{I�G]8"��N&, ֓H��n��\����0s9,����rX��.��mˊH�mX(I�~�)(�V��0�"9�G�-	�os�L����OO�HI�3��m����O��#��T�G����=BM�HGKCC�r�$=#;+������,� �Y�K\ll�R/	����Cxd�E���E�!9z�(--3��9�s��݅�	`88��9�������X@@.)H���#!%#���:r���P|������������(N�Q�<�}��ӅQ�Qx��+��t:V���>>J}�43��<���%$��ed�����]S����70426�������wps����������A�����c^��MIMK�����caQqIiYyŗں��Ʀ�ή�޾�c��S�3�s�k��[�;��\�r�^�V.P.Rrr2r�}�HH��O` �8'ByBI���IN�GG��'|>�%���tǵ�������}�$��{�?$���)� @K:! vv��O�͘`¶?M���ΰp��M�s[olm_C>
\��2�9�D�>/�xY�H�̍����X)�9/�k(��f��UWk�b�V#fFc�[��:=w;�o�M`A���t��t�i��"���mϻ3���;d_}�������V��v��c�?6Ls�=���u��_<���so�ÆP�&zq.��3\]ߙ*S1z+abO�3Kk��3�f9
&f��DCgc'�)Y���ms�]��>:*s�Gs�����8�o'���d,#~z���܉�Pr�@��[n���+�l:�N�/�);����_dvQ?c��&�:-&E�.�w��G���8'�������D� A���m�7��{�l�������4vO	������~�]�yh���Tѻ�!�8�<T�'�r�E�	��S�<'���?' �6ڞ.��<Ծ�I���31�)/>�ݫ�m�"6�����qf�tXxUzu�#�-x��hH����nO�Ooԕ(&>�o�>���?M,�?�z&��q���T��i�.v:ۭ���g��_2+��[�ڮ<�(�����z��nOg�� ����i�ar�`���w��7����#|�r�Rf���Jjfو�KD����N��D��@�k�|����uN��?]:�:"?D1@�����ԥ��v���mW���T��۱8	1��W��
�n ������n���MЙ�Y����[�Y��%!�co����_��e��,x�'�E؅��HgJyaqI��jaƍR�q=W4������[�Ͽ�YA6�6��>�c�vYm��������(��Z�K?�����6`�G�ox6���.-(N:/��p;>��X��z7�Gt�&���@֘n5����J��I�3�C����~�h<��SgN��j���P�3&~��f�?��(d[�q��u�Q�P�eŹ�cQR�7�r%޲�����D(vxj;~m����/�ܶػ__�pض8�LZ�1Kl[��v���&�IXɘ�d�M�a�N)�"aQ�4,����qj�m��.�Oڭ���~'�ɒ��(cY峐3E���]�W"�z�۾$��~�4M^eٙ.ED��P�l1Ejŭ���G�w�ۊcJ�+�{��1��-�vbt�d{���Ȥ�p:9R�>y�呼u�jA���YJ�e���:?D���Sҟm,��U�	H�Ten6��v�K~�ޞ��c�A��"G<�6�U��Bo�#�p�'��D�f�Б������C�D`�ZdO%K�����@�;j8N�|��������-�<Q���B�W��_���i�c���S4�-�D�A7[PO��i=����������5����p�gD�WewH�aI>����I(C���_��'o��=t�gs+ϻ�㚵���#�O�OǇa�g����C�4��Pu��'LI��؊Y��f���o<���w�Qx6�(��$w3�`n����5ak�T�۲v�޺}cK�p����h.�.�����Q���u�U�6Ȼ��B6�-���p��/���-pls�F�ٯ?������z�e�2�mp�$#�<�F�� t�R�_a��{����Fʎ��Cׅт*D~a� ��l9���
f!$c�e�1f��V�B=�q�/���=['�H�CS�ve�oNε^w�����M~�E�[�}B�L�g�dQ\�0�T�D F�p�)�F���ދ���Y�qA�q�P���=���!F@h8-�B��������t�,�W�<����~:��;	�><�Q�}H�����dˣ�@PX���3��&�AP�D���#w-�&��i�0�']�@�x���㱑����%�0�N��2xٓ��A���E?iׁ��5�G�ڮ�{n*�i�?Fo�T�iy��s�R��z�,��9FE�px)�H&*cu^z�n&d���� ~��g!��Oڷ+k(��,�f}����V�#��<��y�2i@e2H@?u�'04�COw�7pپ���� ϧ��1X�ĝ����	d���-Ț)AMh���@�D?ݐ��5pa5��	�ҙ�������4��[ܿL��/4p-�����Ž��I�Zrx^��0P w�W@n/jj���Xa� �*h���?��;�stO�D>f����
�C�L(?A�?ПoS��]62�3|�ō齛��R���ze̷�L���S���G��s�r{��KA]q�W0��w��b������O��w\&��k ����@Cwp�20k�Kb���_�����$����Vy:�a+���<`�o�Z�������U0 ���b:���I������nJ�x .���L��c�#_�	�����ǂ?{��ܤ�Ea��,^����e��ȯ0l|�i�M��]C��[}N-:����c�	:>ڞ�X�ߺ���P��{��[I"���
�"�	. �=��~ڂ�U«p	��o�?%���u�m.2j37bw��	�-/X==�݆䉀V�Dq?p���p<�_��cY���UV"�8��o��w>�O�)�n��=ʀ$��_��@Y��AV��G6b6�_Բ��U��[�
QT8n�R<�5���)~7QS`s�#�(� E������/�����=�}�{ }��+�7y���8޲�?�P��L����Š����G1�D�+gd�:eb��r��6q޹*��l��˻:�*(�
2T�t>�ތz:H��˘RmB����u/нƏ�z�����$��Ѝ�Ĩ3��@�;.������_�$��Z�9e?rf�'	�X-��� �����`�V��݁�<�c��n��J�B?�LT��Q�#�i�\���9�
���%=H�E%�H=[��eř�>�Zsn�d�
WKC�l�|����J��j�h��3*W��-��"Exp�x_uliQ��8&�xџ8o)O{ˎ�;	�o��#L���GO�m?l	>�����xu#~�n���X��^~I��io+j�i����ݑCO���m�������)�7�K�J�����Az �d^?P�O���e`��pt���zK�2]����`��L�{�z9�	��
��.���x�)�?�(՞�%\���#����;����.�V��`bb��g��`kUH�|�'Sjb���cC�f��h��R�9Q+3>���O�v�F��3�#�� u���������q6;��P%9By�~p�����*K�W�ښF�h�K�����g���t#n6��w)�r�c�f˫���s����"Q�U�!�O�В����G��zF똳Č�@��Y=Y"c�#Y.�/ƭ`������*m�z�~|�w�G'�L A=��}c�J�p���q?`�V#�vz���'uGK���<T��S�1}}[F�r�ڂ	���u�J��с�}�|��|��^��!�-�E��Df��ݝe���	޶r�c-h��(�u�YHDPX��z9߶DX���cmkO�g��s��J��P��gek;�k>�ֺ>7�,}�2V<PE:jy/Y/GgGk��g���s��R�<X]��wq*ʻZ���\U�m�R��������tr���� g�y�s��%pύ��Z�Y��;��;�;�߾}���]�����J�涍�++	�;�ŬDD�nܶ���������;������*@<p�����mw'W='�����o������u���?��H�����������_͓�'��u���8�����!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!�!��\��mX߳R��U<x�)��7X��o�#�Or�����<BKMKKCMCCw��q�c�hh��:�p�������4�)F��L�ϟ!i�)�RPe���c��.ϟ!9N�JF�y�����?��M	�%���`8^���쩤/�@�m��u��sO*�na�2�*�i޼�Xt�$��cQ�q"�����Wg;2*m<V7�����ss+]?������l�q�3��]-���{�375�]�~*S�Rvy?_��1���]��K�Z�1FR*�������{�0�z�S�����ػ�>Tz�W>���B8��F���%�[$S�ف
�ܽ'>�QR��U��3)�S8�3���ɢ۽���C-p������p|��,�c�%���i� �k]�<M\���xEZ*�	�^`��/���މ�)��U�.��b	���8�(˵�|�p����<��m���F�!�{��W�l��L�qy��*���E�BЫc��^��%����u+X6�J�p�7�k=�I^f�]��Y��UE����'5���9�|ba��-C�r'U�~�D7�������v��v7�ej:l�#��}x�ԥk��O3m�s���|{�wq�c�� tK6�&��Zbm�#\���� ���#��h�^*1�ݔ����;���L�7��wO�{9�MZp�Y��J�+�QG$�{�����^o�.6Qm>���Я�]$�\B�V�O����X3D�p^������I�ƔK%���3%�\��|�*Ԑ��=�U�؉X߸*u\^�*E�36�k$A��G�2@o�@�f&���VS��L�d���૥����֞ݿD�h�K��7}��{A��h���m�q)�QGhH�|b�1��V�f��D��SV���zb	z��(Ǣ6XT)��؝�$��<�f4�y������O�8r6,�}�GB��
;�z� ��̒�����@+���1��jf���3� ��˝�?+��*V��=$z���ޖ�e��9��vϵ,�L���P�D`,�Yv�_D��մ���_k���yP�HaL���nЌK=�
U�R�wչ���s�����M��QM��1oL�j�ZaaMX�v�2�]����g����e�G�G20ʣГ�Y�ǇX#8�J�&���<�����e2O��ȗּ۬ܖ�J���j��#� ���	<C9t%C�<�z�z<ylA@�z��N�2�%Ѳ��	e3T%��A��8�kni����ѷQM�GyR_ wq.�F�]��?�k�x�Zcz/�ȯg���ۍF��S��b������o�w�֜%M�D�*q���e�ώqs�(�K���2���7<:�l�tz�nh����2��T[L�P��ڍ;Wn?�Tt�3�y� ��n6�|��j��V&s��T-���t��x�ON�krC�B��ǳ��t�G�����yYf��9��m"S2�q�d�n1��Pz�ӳ���Gm�&�]p�te����z���1L�jm�-VD��fN�tæ�T�BB;B��w�av��)w�x{�q�F��$�g�l0�����MݳT$��2�V�,���E�.�B2�~:��In�g�ڱ��&�|���m+-,ږ[I�[��h|���ϭ��.6�֠>��r.���׶�Z�����}V"ИO�e[�s�[.��n��4��h�بǛ�v�؋��rUD�SlY�B�l`��G�é���T��B��Lٓ�{�Z��7�Bl�&�㯜$?�|��,�E�F��EAO�T��WyC���}�:�}��t�����F톧��m��Z�^,<IVT1��}:=���Ŧ�\~-���_���C�}y&ڟt��a��/b�6��;�����}��هC�C��c�sF���Y'�>�Vb�H��-��E>9J }��ӽ��x�F�������e_�p�n	�#A��׫U����M�y�	��;�>��^{O(�s��Sg( ��DgQ�2g���\����'K�r0*" �:rj�M��-ٮ-?5���9�A�R�����}��v�h��Uo��2^�����rz��qߜN�N�� ��=ἍF$�������N�B`R�۫�Ao)-�F���K�W��2��8Y�^Y��}G����'x�?�C�;<45�\�U\�F�R�T0����M���jM9�>�~��� tGv$�"=�xl���0&���c\c�N6{L�9�>i_C���Ξ�Ѵ��$�bm�J�%��(3�{-O3
����t�����L��;^D�:ċN���|�8c�)C8�d�E���Q?��GQ����\���4�����Nu��ZH�P[io]T���b���i�.C��|�x+�i�zd*�!�CR���xP�������k�;�(���Թ��'�74W��$���:΋�4_�Z��ƿ*�nk�f���?������N��	�z��q�}�0�ŒT��]QK�v��d��K����\����H?�ă�[�v8��g�(??>K?m���L�$��g�pQ#�+�����]OiH�^�~N[߶�g�Ψ�b��Bc̛$_�U��ny�E.N��iEޜ��lL�<���r��1h���Z��Mӂ��bI��/�I�b�E�c�W� _$��oGf���M�r�J�u����g�׈bG���A�!��|9+:�	�l��-�^��h7����)������_ݷh��P�� �Z^�=挹���ʳa�	on˧*g���'��	�����؛�Y�1�4">���Y�H��N�qP}_����������,c,E_����[cKFУh�x�'�lQ_��I紀�5��BC:�"k)ŕʧ6��o����L�Ό�X^*�M�=_j��v���$ɱ���Y�ř�g(��£b�)��tr�ڛ����z�U�=o��=e�V�wS�o���i�0��-�����y�V�ό=�}��ղ �Z����Ci���?ӬȼIZ_W�����d�E�BZ�dH�8��vΘu:ۑ�~�~T�E]Z�#xX6j+�۝�VT~�/A��2���������G�5��YJ�a׬�ʩ:af��ى��O��\-?�q�z�8_|̦K�м"�zN�R�ʋk���Z��1��*�[�r�9�0�U`7��+֡����ɡ�,�A,i��n����O����8n��v��x�[�vq�؍G73o�_ ��u�&s��k�9�,5r��|�K\�=�A����'��-�u��I���'F�9��޲L�*?a�Fl����B`r"�̈́5�J�/t֒6ۃ���z�7gY�tsZ��[��3�}��W��-�ؽ�ǋhX��q5N}�S?v¹��g4G���3���!��Z��YCj���*'c�?q<�Ͻ
LF ��K�Rk&��G�x,zq�'��aa�O_�4HK\���_c���A?�ӥ�\���IT[IFض;֤�#ͥ_�`��}Ć��J�#�>��Nl;��3풫R���v_Jh��9$��Z*8������7�
#`;q#8��:oǡ�-�b[����Ӆ��V[�7�*ո�D?�=���YрIϓH� �<���D,x����v~,6U2��%��1�mc���@�d{���9.ˀ��3���޻53�%�k+1f�$C�o�}SxPw���8�z��m.�t����>��Cƭ�SY晑�a�YS�Q麃2��f�s|U{�^\(v���)Llu���E��)��Ky�Зe/��kONgӈ�ce��yN���Bf�9ĸ�i��*o�!�n{Z���W����\ ��Y¿���ڥ��*����`�1_u��ޛ�r�{��=���[8|���S����[}�+�[�eF�S��E+�(+�P��S�o�3���t���]�ԓvIz.�kΠ��El.�s����SK����N��tRE���Ӈ����
^�0�ܣ���ѹ�	g��n,�XN�\���I
1��~���m:�٢�\`2ӕ`���=�c+�2^�|�Ơ/��(��x��5�<"`�g�n@��X���.�Qo�A�flN^[��xX���Y�:ڣi��Mi��<��e��AAn{��R�R]������D���O�f���H���L���@��@�3c��y(��s_�L̛ȥޠc��!f��&)��n�~�rSK���mf.;��e�L���g��j0��?^K�R�=�f<״���լ}Y��/�4�������\V�:s�J�����q�'�ߏ�-��32�1�����H��Y1�Bd7����i�DM��8���W���c��2;����q��F������ꑬA��W�i�{Xڢ�D�1�)O]����*.������q�ܝ3NENt�/������&�_���7&X�g6�����Ju���:5�]Zn<4� �[(X���\]?2���c�$c�l��V݂G�z����c����q�"P�?|-]wY5�Z�X\��D�v!ˋ57�s�t�;VN�w[��,���Sf���\��/���E��)o6�@���0��p����7% �7%�/~<�����/��S�ԝB%F���B2��rҢS�x~�D�P�$�+�}j�<c�7��hy56:�������}�D�K�N��R�C+G2�T�c��H��=�m����s��E�W8Y�Y^e�d�þ�pT&Zn^�M�$[�s)�x���7
���R��4�[��y����R�����(��5b����O���V���^�p�~��M<�/��薈���r�UԴ����SV��5hP��v��;�P
��.��i�C�t�s�FU����(>W�WE]�,��(ޑ���^KĘ���sD`�5�O���U�����s���M��h9�(ljz���\K�ƽ�m<bcπ�L��{"�G��L���ct������,���EB+u*�-޼%�?Sh�D>���+d|��-k�Jŵ��|��?��̀�~���x�f;5BQ��
�D\�a c`K"��$Bn%(��D��B/��M�\ ��e���a����:qF]wj6$o6E����E2T�8��)??��|8֟�s�)
EGV4�^�6O�D/eԐ�i��������ї����­�	����{g���7�nvO�m��D��w��1�}d���%�+���v�?�/�ElV��W�H��XtՏ>�o"�p��q�w=�&�d}��SO���i7�X�7�d�F������KD ��������Ih�L�k��Lw���I�5��J�� ��_g�ޞ�W��D ��0��$�`��Z1[���'7\�]�� �C�WX�Z(�'�D؁V��!��X����CKs�3�i���Z���M ��U�v�YV3Ia���i��#�(uf.���Q&h"@Ͻ��M %_����_�?�A�E���'w"��BL�QEбI!��/z"p�ƊV��G��g�Z��/)̴ߕ��|as�S������grA/��>1�!{��D�:������M���s�-
j���1��ضG8��]�H@˪�xb �B8R(Χ�'K�h��o��=1*"��;�����w72E��
��ɭ``�Й8��ق�&�!ۍЫG����(����:_�|-Fn,�����@k G����'��~���B��k�����T#n4
���yT��s�����G�Ml�����`4Up�9�������]q��"=ƹ���DZ8��2d��-��(��(�7�����ӄ��uk_8���VK`D:#۝p�`���׈,�\��g
��:�4�oF�p<�D`���{�do��l��#A�l^��=���س}o�]2�M�L�S�[�B�s�+�/�[ٳ2�J��Lc迕QO��\nK]:�"o���p:��p��p�D���Zg�:���u����1�B�H7I�I�.�K��%j.	@�X�:�����~�\�W��ͨ�����7	BD Y��F��֐�SGK%;������G�W��fy8�b���G"�ǉ��h�<���q�_�tm%]d����[��aϪ�p/����JkL�x?�6�{���w�ˌ��ar��k��z�����:
�n��ې5���2x�m�	~�-�����q\1�J��܃���5����(�G���7������Am�ުe�or��㛳-u̓k\���f�|ߦ��*(�f|���.�-I!��DyO�F�S�����S�)����_�y�U���y�����Y���F�.|��eӕ�ݢ�k�G ��Zw��\u�Ĵ�1�KԘ%b�[��P�+$����[�S�Q��0����L��;�H�k��ص=��[�] �ź�"���3�\oN~&u��l�p�G�����1+
���RzW��������v�����c_�^�,<w�c[1���S���i��a'Au��)�����a�����ga��@q�r�r�GӴ۽��I��҃��i޽W�]�����^v��idw��N.i�����Q�Q%�Ҿ�8��Њ$�EH�ؗ|��m!!����T�J�Ov�4=��{FI�h=�a�pv4:|Mo*Ȭ@}����N�+��f��|&��2���{}/�������Pn|u&��#gQ�����d���?��+�O�L~(�7a�u~f���o��R�O�;���S�����K��Ֆ|YЍ���]i��Aгa���/	���Yaͅ[�'U4Ce�춚�:����a��۠�YA���'�z)�Gp���xtB폚>����ox�h��/�Gv0 =�Ϫ^�C0��"���� �#�I��D�HI CH��/��C�C��ߡ��pv��J
���.��~~b���a(���B���>"��³mM݊�����q���H��������3j�e���[����G���B��'�ye��cV4��s&>UzɬXR+���+��r�^�[t�<��ۚ���~��M�����+����^;.��G}�i�% 50R:���W���$�^E�x~H=B[�x���4���`9S���h����Ѻ7��$������V����k�Fu��*I���Z{e��*6�!�b���zr�8�_hImp����O�i���N��*�o0|�'��s�:g�Ħ]��qבʖ�'��e,���X���7;bdxkn���>��~����I%�&��%�4>���\;����}u��q9�5�ڑ�Ua����v��Q���YL�i�3$����i+v��fI\��O6{�u�������4��j*���Z%���zQl���M�(�c�]jU�`�Y�������s�l���q/������&�f{>��L~��ēouu�)����i]kr�#����9��A|Y��`�1ѹ
9��u�U(_%�w��-_Q9�Ys~��J�B,ǐ�7	�b�;����|<� z%x/�� �C�M!5*�� {���i��Edn;�/��e�}!�\���7���ޯ�(�բD����������0��_d;��!ԯ�?���LJ�S��o~ u�o�߼&�8�O���	��x)$QHO��/e�����Ω�}}��|~��H��Ek��{SR�g����=(��\�א��Or����HOc�֮�W^�Ό6A��;|=��u��q:}y�U�&�-d]�~v��ƺ>��R4�'�}#f��T�
1�ml�]u����Ϊ��H�\B�v�w+Yt�B��;c�����E�u'����-��1Ŋ�`���Һ-�1���E���v"Ք��C`���^B�n�1��Tk:��2M�3jՓ�?I'�ڋ}���1��܉��{�Z����슗O�c�Cڅ�C�X�7ܚ�V�F2��>����h�m�b��er�&T[� �o��{ď���y.�ȉ�r׸�n
��ݙZT K4��r��a�h)����g�.+(_m��~����쨁z�Ԯ�_���st4iъ��Do�Cz�
���xO��Fka��_c��>�h����ʽk�Վ.���`�0*�Xi�a���\&3n��D�c$�j����a����8Eb�t���l���7O�͋<�+�%��B��`�)5�0�[\{Vs�������g_v;ܗuJJ���ؔ�^d�������Hj�}�G�h4��v�b׹�9.`x�kEk���}��	7 ���"�3ߚA���0��H���;�<�|�i x��Z-@k؁�7�&d�M͚�a߸N�����kj0F�p������	�ٟD��ϿH��N�I���b�.��n��quͦ�^�Q��UTG�	��~��ᴍ�����)��Ͽ�[�g欌���T�6_B�"��R{�(Ȁ(�j7}i(>o���$�O���k�6��E)�񂪧��r�."�2	�1�Ė��&&m%5�ƒ�e�%No�B/���hX�`��R�a-*N<���t2�2N79X(끌kwT>]dA����9��$)㙢.$�U���<��r��M��?�|�����z��� RC!�!UŊ��؇�sn�GC�W/o�D���om��h���F���;o��\[?.e~�r-l7|@���~�?�@��P�X�m�}A�]�.�M�\O������_�68��/�XuN�B|_#���?$��|�x]$����7S�i
��ۖх�����D@#d^g&��/��(�=X�O���F=�9~B?jq�C�Δ_6��mi�]�Nl�3�25:���x�9s/~#�|�M�ayث��B���8=lW�4�M4�r#c�ߨ#�#����:��\I�y_C�|"[_ݚ|��jj�9��`m�K�Q�e"�`��
�@P�֜E6m���!#	<U ��1�2�;����JppB�=�[_���{���N�R�]��Z�5l�Y"����Pa4lK�ʨ}+���"�Z�C����B0]��¥-r����D�z�u^��G���V�A3�3O�eD`Bߡq��~�6b�VL%4� �RIUFyɰ^/T��&|�s=�=.Y��|��05>m|�����{��rl�?���Hw��h`W��}Zg� ��<�C�g�y߰gX^~)m���o���?QŮ�jk�Zl���9�>
�����*>sC;ҙ�^R�䷺�S��x���^��^S	[�S\�H�D��E�����o� D�w{\���~��G�;�J�"�ED��!F�����n���y�m��+�K͹U�`��_�w&�˯q�1~d{)U$��;gX:�xZ�W�U<��{�0ɭ�HWL�Ub\S�&��=w��v����ocw�n�,���g���2��)c������!mM�t���g���OgŨ��BKK�q��ǡ�!q͟�]���G�����Ƙ��a��n�X�е[TϦ}���6x���2Х�7v��+)]C>�@2z�˵3{9..���D�^L}��|:]QV�y�Mџl�N��c�7�ǽh����wm*�TPZ�6��zl���	&+2�Ǔ����]�D��k�c��;��l�h��q	x�؃��|�{p��{�=fY��w(�D6v -نV��Z�/�[nD�\�>���|�`��d�N��N�UU�} ����Ռ�z/ [D`�$�}�Q	D�ڒ�9�i���
�|�� )��$�+�u/����iO��s�p�{S8�?��,�� ���N#"�{=�.��.��N�2�Aa�w��=I���S���LG0�H�vf�
u�A��(dy��i�hX^R�v J��j�@�²b ����(�FUD����of�	��$_�D�%n}e(�[G�I����¨Eb�2�	m��	"݃x���I�*L0K" ��#ӯ�xu�B׶ }�z;��Pr#'�:|��fӁ�h����͗��-0ì�Ƌ&����aH[�*Yzb���3�l�C��?�@a� ?��k�̀l|K��vIn�#1��1�3b�I���
����.%�E.��}l����~@<�¡L{���ߍ ;v>\��/����jY�z;#�*�k�I��\ne99��<�4ώ��}���n|�w
wK	]����nU�XLi�Pz	5oJU���_����T[h����	H	�=L"N��Z�⺡+��5���T&PT�1�� Tgw9c
�%�:��EF� �� �B�,�&/��_���|�$1{h�j�q�47��u��C����h�id���<�jWԐ��F��qN�OQ(�}[.���Ӻtb/Ț���
�"���j�ɐ�,�M���ֆ���7��?'\�1;�t�G���&�n" ���L�?�	�C?f�ݑT� � +�����I����j�N���F��/S y�0`@_7���#ς���2�_���Q>u�/���gL	搂F�x���ǜ�x�c�l(p��'�����D�'%�	
���i��P@x��������N����w���@.dl&o��b��#��絾�����H�|�s��D���'��t�pq��#����'�Dʋ�O!�a����L�$FnI��`L��@'��ߩ7�U�N���H��V鰄
秶E�����~����I�g�l�FO4#GQ���1"`٫�v]�<~7�i!�@P<O����p�����LS@�9z���ǧ�4λ}����R����)ws/{3�/�>%��w��/�A-�r�4���ܕ�u��i�K�T�@%�y �Z��xq1%��7�n%޺=J��9�\"�ĺ���F?�5*��V|� �}3�U�fsQiaM�O �}G]~�Sdݤ
	�1�/7^��/��L"z�+��=�bDUH�(*k]^��N��d4�����W�4�J�����c���:om1��n.��[���9���E��x*f��׸�/]-.��*�ᣂ"/�m'Ew���l��]p������n��]���	�H/�M�x|0���Ʒ���2�X{��9�(�c�ȓ�󽋹�1��[�ƙ��q�P�6��O�4Hp�57�X8~�&@(6luZ��v�\�Rێ+����0MbٖA��i���[�$�vLK��H{⋲$5�K�k�Ü���{��_�d�7lA�d���;�?x큼��I=���q5mq�}��"���'�(ԏ�3��j�i�,�7nn�_�%�s�.��W5�p�����Tk�.B�кG��\u��o��m8��\�I��;��>��*�2��]��V�3�=����e0�U������P [tC�K��f�����h���~a�3�G��R:"��Q���2W������՛b���a���/�]�֙��F<Ǯ1���_�i �?�&��us,��Q��^%~��p�}�t��(g�	ϑ��kg��UE��q웢Ӕ�w3������|���	�^����V�������
)��͋�s�D.��=t���Ft��"��������|����G�s�gd>"=�.\���$۟q��6� �k���W�J�_��E�e���b(���=WxSӐ�#׎thu��ƾ"�eA�3��zD)G�&���;^59�E�_-''|��8*���f��L.�k:�Z��VV���p�&��N���|�d������c��[Ԋ�&I�g��H��n�D��Agn�ދ���/T\��``=�MG�C'}z���9��ǟ�@�rG�?�]����F�RV+V�~&�"�xS"pYbnkrR��Ʌ~�����Z�~�a
Qg����:!�A�6�d� 4ЁY��U~�g����[ݹ[���ȶ����g7��s�\� ��b�
���fƇh��L	^�=/��k+ք�93����ll���W�w�5	3'���7�?(2�&���i��޿tMye��92ҟ��HY��9�{Z��LPL\%�Tr��<�1!ى��|dO;aJRLc/S�����C���`s����������S�j�`��o���������L�8_�� �9��Wtg?��:��vwc�i,�?���X!��Ad؜�&P/|�1��}�ę�h/�R��vI3�AG�S���S�K?�?_][qل�e/����	���W�0��iA]`�3	�� ��NgI
ޔ����8d2x����Ff��C��e6�f���;���LIP�tg�S�����*������"�ƃy�)n��?�Wd�a��+����'�lׁ/���YL��k3�0w�������p&�����oz�N����t����o4v�Y�����f�줫_�f~=�$���=h���]���,Ź]��� ��Ura��������j��o)�І*��0��I�9$Db�'�4��:쬺ͼz#$�-j��Zc�����_T�8���-j쑍�p��Y�������Cc���=�fɿK7��E��?�a^��/�yU��-dUhF?��&4(�Z[���qz�[�5ݿ�kk�ħ��u��j����6R�U��+8_���yr�WEQ�����l��Լ���w��6�ֈ@Y���^�>�W���l�e`���/s�$
�/��;�t�>׬G����#����wE�77�*�߮i��	���L�俥��`J��!d+��G�k
��!x��O�_����d3H���-���`����Z����c9�Q9C��>@��o��B��Q�-�a��D`�$��ձE�X�A�Wg5�D΀e��ڹh�־�K���╢�T*�rf^u�P	e*��k�.n1��J͉�-%L�K�����ڸ��0�q7��\���ttB�{�w�w}�Z�Z֚Y�5��y~�������������_��լR��/�H�L��g�M�v�߅(�}���ͻP˿{8�\��S?:|`/��H}��틦;udL��QZEXLVy����sF�����PV�Q�
��`�p}~PA�@��zs~�a���;���s���\7QB
В��·K�%��6m��J��NFiO���y
<̈�!����wߑ3���Rv�w]V-V���'�P9�]��PL�������H�����W%��H6� ��.��"@�<tl��u-�����~Ƽ�u/�^
�|�qM�*�5��a�\�_�Yx�ݸ�ݪ�7`%�1C��I1Z�v�G"�))�*dז�Lj"�"�T�~�-�s��E�gD�_�O��{�����6�1�ܾ�u�7�}3>7���m��<�/{S4������*i����ѱߦ��d�Lg6M>lo+��-"Ç�t������X5���+r\���ߦ��;�{�|��]o�:����U���O%��ȱ�3�&L�<M1L�ml� �/���V��o���A�n7��?���V.7�4���d�w�s��u֓WH��I
sy�n�Ks���y4�u�?TO�[��ʞ�p=��r�W=�Wr����C�I�6��tD��ؓ?\�C��za:�u�@�ewoPD.�^��eS�}ɶ�#I�L�>#�C���MpJ�5fpxDI{�z��j���1�:�B R;���t�O�@�3�=Y�փ'�A�J�>���9Z�N������u�ǺH�А,����`�9"�2���SX�ѭ�bR����&�MYB���`�e������k-
��F�r��e=J�7I�s����P�UR�޽JA�0���'ꇆ�a{)0p� \�ۆl�/�@�,���}O�{6���A��%\f�vv
nL���%����ڽ�:�,i�P�xW<g^�����ymB����=�<b#�'�~A��Eg�p(D|f{b�KG]E�"��x4xO����v*�E�2��b��w�%0��%Too{���(��f��"�N���ö�'�"qw�h�5D�_X�K��ѡ�QȾ� ����C����/�������_�G	�k����^7��4&�P;#T;�(��qAe"h\!ՙT��fFG˧XBj.:��w��4,��GD�#g�>M�a�T����Gݭ�r��leHc"�	���	���wZ�i����W;!��� +K�G3V,n�U�Mk�N�!���I��3I�G��/����ft'E�{k�ѭc��cu��Ƒ�1��.�U��[Ɨ��
c[�����u�8��/�@>/j��z2�	�$��������Z��_�|���!U5;�)^����#U���`�1X��Ar
a=�6d� N��&4��wk���4���S�툳����*_�J�B#��廷d�?T����������~6�>�p�+�H#�j���ay655<���`���ux�0-�B�D��s��hC�p.v���Tf��ĵ{&\�G	G�|�3�r%d� h
�� ݛ'�&�{%t�T�8�,KI��j��������q�HNw>��t�ӝOw��w�b߫�ds�����,Co�I �;�jj��n� �C���;3~��lA47�Ë����b``�N�3f�UX��r��kqXץ8c�d8�xi�6״�A����&=���U���9Y�/em1��c��R�>�-h]����y��
Be����W6�%_`](���P�@�S�`���OF*T�8�����˲�CH=1�7A#���!C�\�f�\��s�+\�|�i^?]��7H��8(cP�o�!o3���'�hN�K�Ӹ�z�O��HI�=F�j�l��~יs�`U���Y*K�(�F`�5�Mh���*gQ�_��qW�a �M �e�[QA#��)�r��d\�ַ��2ED[�����a%�%�Vl����j�:m��jS;-�*`�-y�as�~�I�)����n�X[;R+uÈ�T�1���G��t�;��H�}B��<��ɯX'����z~���`@$�����C�-���(�P��&D�!5���bǡ��x$��h�*�#V�ED)��	�]�&�����g�U`�����a��r�XC8pJ�DQ�Mk}e�˲�����:v�\���3��d1O`�\���k��MJ_�a�h�$O��)��OM�t*�$��
)���H9IS�i��c�R)󪫟d�D$�\��K?,�T͔Pc��T赨Ƶ�~Dn�/żYK�ݠ>�S0*��s��V0P�M�b=/O+^Lk �P1��W�	tA,���;�ū�a i8l'��9�c����R�>nx��^BM|���N����/V�6����0�p��K�ُ���Xtv]���;��nr~J�쵔��Ӡ�>��ײ�����}c�Ð�.��T"\��='�]��_JOr�``rp�l����]xvR���It�����ɏ�v��h�Y(�6j=9s	!�I��E>�m�	��<Fz��~�G�_�)�	q B�eK�j0����h��_S'������}'��?Z�˖h',f�\�A+�����=|`��6E�.ƥ�o�`�=�{����T}��U����[0!��"��OV�7�X��0�f�関9�����܏8��|dN�&	(�������O�qЀ4*�x0���h �u	�"��j��t��[|����od������|VGU٨�T���{~ {�u90��.�s=0��L��c>u�����Ñ�P�Gi��U��T�#{�F���͊>���.']'s_��?��,�,i��y���R�L�	#_c ��E�q�M����;/�}����3�ˍp��Ga�;�2S�������V�9��A��X��,�#/�ݐ��z[v�e��f�����v�꾫���U��Ϙ]�M0���,��s.�Ȭ��`˳�s�N�Ե捩7!����9��r�����-`��'�Wd��7���v&�Ztqmr�;kSy�:v��X-�/��M�c����L���L\���Z�)�D	���g>g�[��q흙�F�$��"#KhG��QD��U�$a)K�jP}|q`։�m������nTUʹ1]��8o�0(߲ǧKYч�GyY�|�7�����+i7��rc:���+����\����aM޷ӻL*�hq��WV\�*����G	��{l�7�q*�R��j��N|���R����'�л������r=�Oo�z�F�E�s���7xt$��G����ú��:�d�z7����>u(c\P�_>�|��%7e�i�]]^��w��"��W�86.s��~p�����,�qύ>3�Q��?��+��dӖj,��/���M�5�R���3yL��0ct�N����F&�����ҫ���U��?]���tYg�B�g��(�}��7���nb� ٜ`����YnMF����au2h-��ʕI�x]�z8���{1��x��Q�G+K�-������K����#e�4a���?���j~o����fp���\�:\�Q��-,2��_��2?�;��Q��c��Ö%�%Nkb�<[���NY�N*��9X9�����nJm�
V�8ET;�Sk�;ԃa$���Ԅt�
�H���wo!����
��ފۖI�9�D��H�e_��3��w�沇����`�,2�R�����F���*�������	FY;���i@���qR�����I����9�"��x�P�O�#a�ꤻfoCR�?�6lC]��fZ�(S;p�����~�䲛�k�S��!\�5�4�i��������Xc);�,�c�5�բF�^l'��PE�xR�)�x�5�>S��<~}��3�zũ��]��<�8
'$Ӆ��P����X�����Î��s�Iw�i�ҍɼ�[#y�8)�w�4�e7R�4������j9�V�VO�o�o��97Uss�]ME�k~j���C����ԟ�,��-򊏂E}|�'+ؚ{z8���kHvx������̝�
�,߯���`V}��o�>���\�x�f���n�s��O�F<A-d��� sHg����+�kx�h���PK   9A'UD5�<� � /   images/bf05f532-b4f9-4ebd-a877-7859e21a15d5.png .@ѿ�PNG

   IHDR  �   �   ���	   sRGB ���   gAMA  ���a   	pHYs  �  ��o�d  ��IDATx^��dIq��U�������Yo�u��#!�G q�8�� ��;Iwȝt�	�I��'�@�;�.^x��zo��tO��������W���{zfgp�љ/322222ҼW��v�@��-Xwc�*�.��鶅�벆>�V�/�������ln^i��銲 ��o����#-CW�r�Y<�/*���T�iSZ��r�3? �/�?�.�G{z��O��k�e�gaQm_h���ʲD���PJ�B�	��"O��UU	�%��JB��2�P
F� �V�H#�\9�Y��8��Z@q�R���ыh�h�b�.��7�6����tuU�)�e�f9A�3�YO���V4D�ʺ"9='�8e�3 v��%p~��C[��Cl%�C���!7���6���]�[P<r:�.���%zz� ,�
t ����w>�W�x�_�lq��Ҁ�(%�=8�r=�+mY���HR�Jo�.Z[�r���9����w�B�Q�]�a-@�3-zU��&�]��V��)CHw�A���ܩ�D������v�P_�Xo�-O���ذ���d~_�ϒ�V��|���7���yi���y����k�F������92jS3��b��n�|�tƢ��ieh�<h\<:���N���E��'��CY��O9�4�Ӆ\��0N�CƊ�06`9�R6����*v'����03�Za�ݩ4ޝGn� ����|(C�CzK��u�t�e8�p��/Ģ��-NITK�ʉ7����n$��Սb0�I���bGŗ��Qƅ�,�W-����*9�qP�Id��ת�\�S)��!��,E^���Z\ƠͶLV*K��B�p.�С�'�K�C�N�v�Z��&����k\�2%X��}�J���]��p��c�j��'?�$��8u�oUJ7i�N��:�H��|���,ZH�e� %S��	P1�	���I�%yy���Y���ˢ�I^��F�	��@9�}��m����>.ңl�`��~)[���X�+$ZS�f��@z�V^��-�=ds�ט�Z�[o��6����������Q���cvm�3��[�ѩ
���3��۱2��\)rA��2�{���)�꽇��7�n_����N��_I�*�B �>�(x!\ģf�zQb�9L�ţ��1ez�����Pl۠+AGn��S���U��B-��)�$���a�_'��B�_��j�!j9>-�2:�J=-]�j;�	%C������2`$θ��IJc��@�Bw*�C���x��c�RjAmA���]�%��~3䘧����ٿ�j'���W��*��۟�joQ�8�|�Q|Q24p�����Ot��LsZ�r�V��	i2O�x��sR��1	� 8�z����m8���A��E�Б��>�(��c"�'T��M��L�����s�0B��ԹYU}S�"�I<�1�D����U��RD�3��C{�W������+�j 4���M�=_��IR��c�����)~�2�$f5���T�uՆ=��s�I�f�ܽ�v����O�BÍ\}�&{'8��C&$Zf#���9{�g�l����gf����4[V5[@cs4�ίt�@�$��uy�!�
p��9�s"��x�,�K'XB/@�c�.��v^.m�p�����x �Z΍bQ��uQS�eXN�v�2�Q._�x�������;ʒ�~-B�/��
�E6����<墏B&�3J�1P�ZY���n9��!2�N��>��t��]@<v����+��6$�mǽ-��"��*���|�E�� �_&�	iLx�>� �[�>Q$@�%�����|�OJϻ��M:ta[�-g�I+��nJ�]�z�d��X��R��()���pk(�ߪV�U�bi��}��s���cQ�b��b�P�Sx� �vdhgAUK&a3�)W��M>�x_�;*"ea���/X��m�M�ʨj�8,�3�u�c��`/z�U�km�4(,���x�q��J�s���fju����K���m�b�=�QZ�حU�w�������#HBO��Q�O��24\�ޡI�z��0rr���'ހc@K���u�N|�&���a�+) �-^O�D;��ˆ�x�q)-���j���r�&A��>�|�0r���W���?ڌ��5�Ex9�����NO�]ѷ��bL�nO�M�yr$^>Һ8��bY����0TH�ݎ�!Q蓍�����Ę�K�Ew�VOz�B���z͝r�֐Wt��vp����P�縓:˽���{+GEȬO����Cw~�nC�Qf��`O߹p2,hG?���,N����Ɏ�����ì��baR�z�.�N�V����Z߈ժ�Jb����6��O�RG��&p���d�'ȋ��A�fd�!�V'�)B�'�Ԍj���J�rībY�μ�t�{N�K1&��z=��f����=�f�{�3�	gm����G���:C��G��qi2YX�ڤ4���������Ikh��K6IGǌ�FU�A@ģ��Ci45���ID=Ԉ��������JW�_G����3ӆB�
"<�ؒ:͂�������)��x��%��"�Kn����FeR����Rq��h��w��LNF*e��t��\�w���4��uxN2TO"J�0�c~�t�A��HJ��:� &Z����6U��B����OI�_z̗�K��&p���%�{(Z����2x.I�3 �H��SDAa��d��Nr�>k�c6p�럝p�h��Ё�Q�,����c���p���C�S�4�g��q�VN(���EȾ��0ʃZt�*�~�
>a���ݮ`-�'�!�g�R{2y��ݭ���I}�Q���[\��l�t����j��k���;_(ΑVLx΂�B�I�I=��4�^���E�!�l2�����/����~g��y�ו�.%���OR�ZZK��u梤T�:Z�m��㶽o�^x���+α�����xh&��
�'�lh ..T���Y�������=Gm�n6U���J��q��B��UT	Z_��
iv��Õ�9MHJ+�	�n½�q�R�]܅LP(X�|Z�bd%���$�\:��Ї礐2Y���uF�V~�q'����U���g'�늫�m�v��PN�H�wQ
bn�}��r����9��P4r&�@�(�� =�t�X�[Qx�%'��2���s2A���%�#�<OmB�$ˑf�&d!�ʐ�^��)ʊ1�Q �/�
�fG�2�J���l������[���N�q�uO�M}7�T���>m�2F� ��˛`%�2,�e%H:^n�3	���n_�X(��M�>~YG�Q�����M�;�Q�����mz��U�-)O�e�HQ,,y�j	x�R�R��P.C�)���:	X�h_���誡\O�#;����?��]�ݚ��lP��F�=vO���%Ϸ���R	���N�L>\�i�ך�n�?n���'L��#ʚx���ܑ0-�lT'�!RBx�b.C�w	H�%��[�>�)�G�r���+��^�K�\�/h�-mj��H)H�|��/` ����b(`x��������r��6����������z�JF��#�����k�?<鵦��|�ߴ������*�O��!�,:���J�eG�#�0�n�^����p��4w�4�Dft���//b�KB�(�&����`�m�9b�c�g��,�{;���R(Ȍ:@8��e����������e���>h"��Y�D(�%���O��)��Y�kXQDr��8Ed��-<�O����&b��m�z��¦�ljׅrv�6�ݣz����Ӑa��͇�sO%"��K��Nd: �ޝ�W��:�����&4ӛ�Lȸ��8�h'�X��˶�Ͼ�j�d��Ӛt�Oj�ږL>��ֵÙ�/��_��7�z�Wi��]@��q܀���4@��0�A���f]����c��٤���b[�MU�uN���v�6����������hcP@e��*�'��N<�l+��	#`������Sr|� oh2B!�����F��~'	�b3�d�r�,}�j%��u���h����m x�NV�T��j�g�-�F�q���&�s|t�B�k	�b�E��+�y�kj�� �;x4�t�=*�e=�GV��бh���6M�5��mx�����s�qV�h��5�CH��}OJ��|��{H9����LOj�"�Nd�iB��M��&ʓG����d*���G��y� ���aE�:���b��#V�z�5N�c�6��_T������A2�e��1'�>I�E�!��r^�[N���l�՝?Y	�-y��
��-�{�eg�c\�8bO>o����^`��f|W�}Q]��ɇ(�ϱz�����?�����jR�PI�ėL>	�q*L��j`H���z�`���.�*��r���8+���D���D�b��T����s��	'����?b]�<�#%P2F�0�; h;��� m��6�*n{�C2��M*�6�Q4S��cwn��"c���� �s�2�đ�Iƶ���t�7�K�Q..c�p~J�*��/Q7A�;y���x�-M`$�?�lrY��!Y4QgSF��k��������Q�������z�7S���wY�F��! ¦|J�PL>A�t�o��!~��/M��M@���ɼ	����:W��Z�U�G�]Vi� B�M�y��}��j]� ]q�GѹE�M�:�a�q�Z2-�#-��v�����$s?9�l��-!K����rz[?I/�{P��F�b�9i�f/�Y�W?�6+�۟��z�b�a�h�cs�n��uw�/���vhaX���E.r�SaP��S@�DM'���K�^�S�J�ep�<�D֩|;���"I�}'�v^���#3��フ4:��`�lH�����!�Xs#����t�q�Le��r�ONޝ*Gf�X�|��iĉkg�KL�����N�@�q�!&%"ſB_�}���?���^1m��|����}v����B���+��(φ��ũ:�_��t�F\m$�[��}�k���rY�8M�Y�I���>e1u�5��R��	ʓi�bnX��/�.Xc����i�v럟�9<�y*��n(�ڽ2D��B��v4�D�q���k	�[a%�v�&�r����6���H�y�L>�J\//c��-���7�A���V�;�2�Z+��ݯ��_���Bթ..Á+�|E��b4�'�%��	Z ɾ�q��TvYh����e�с_��ns����nmZ�U[o짞}����s������*u@wY��f7��_|��3�3(#6� We<�]�~OY�( �LMy�Ԟ��P��35���[	��򫀲<�|žTo����ЖpX�>ږQ��꣐�K!4ܳ�a�p�Z�V�ҳ�eC� �Q�W�;5��%�K���9�84��dC2�Z�@�ff�mxd�M��Z�/�+�ʺ�9;��B��n���"�Wʹ9��>�0l1�B$|^S�J��tu��?�*~�l�ԾR��n�ab�h'�:�!��Sm�'k����4emr����H�I�����Rq' ���kj�"O=)�/�����p�b��$�����*��A��	qA+��F�6k�34}Ȇ�i�=�5zչ�|����o��v|�F��_I+d���!�'^%p�U�ح���{ml��6���U���oYXA_4(ڇ����A���/��	�E��Ivu����/�2�o��[�q��k���4��G�u}�k�~�]�q��(�,���n�mV�[������o�qW���b�sB(�U���P��3��7c�ʼ�\�J���L(��D���rf�u83�
ʓO�X�c�b5�N]��B.�a�z4��kFjH�~��l�'��b�'*�4;e�f���U6}�^;::iW=�)�w�~���O��������~��*����$���9��/�#�&�]��Q"��Ӝ�i�%�32@��QZC[�I���6��C�*|m�H2�Va3�Ѯ���ks�����#���Cޘ|"Sa갰씾��)����}��RZd��A϶�C�$[�����q@C����"�ޅ9[3̶N���)M�*���Ǚ���i��� ���Yp���e��^*�j��ɼ�4�7S4���Nk��h��h��~!����K�lH((X+MqoE����|��m������,X����8g}�u{֥��o>�*�'���qYXh,ֵ�Y�{�����~�ݽ8,��
JpV 8<As�1���.�:��N�������X��Q�ꡝw.���Z@�Q�Y␭���������CW��z�ze�$�GawN8�� w|����-ӇmM�&�\����);�8}D���c�I�	���x�M����#���'=����ﲟ��������b��q��ܟC��oI�� ���?��'�h�B&�f�;+oT�;!�Nz�8fj��a��j�6Zy���(�����Ժzl_�f-��|�{����p�%��GJn�����H'"]��BI"U}���虢ᳰP�KO�e�8�zA�E��s��W;�Y�8{�q�6���Oy��ϼ��ܠos8���u�ci%߰j����i����|�UGlv�e6����2:���&�^��#U\��ăCe��ic�-�t�"��	��w翜��*~��W��Nݟ����eo��g؞�#Z��A�uD�&��|�sv�.G�q����Iy-�K�p`tO^Y�%�.��p�4+@�6HIM^Җ�6(�j�0�R��!iQKQ���P�#d���ww���|�T��2�n����S��C:�U�A[;'�?dúvT�����7�����Y��U�q4��GP�F���*6T�Z��T��ğ��Ug�r�|��%Mؐ�4ď�b@B���V�3�e�C���Ux$��nN�����@�[_���=�jc_]������������ͺ�î����ld�0)�q�!�Ϊ�>�Uz7�uRb� �$�75��9:+�ϔFz`L"*�0�V*�������uF�x�c��NG�����4��g���̫��=��>�N|w�� �w�q��gv��O�\'�,w�s|��[��������Yd��&�����똷��ywMRGȅ�A�o���dl�B� �~YJ;(��8S�y9"W�O_�IItri9��P凎�ص7���W9б�䀚�kЅ��1�ˠ��9�\�����.>.�K�I�2g��%#&����G	t,���2D^��;���a�m�&C���+
���q�S������G%($�~�e�v�n##�ln�f���֨ˉvi�P�z��_L<�������z��U��>�&PJ�J ���l��@☙�SRdB�̺vA<��y�V[�mV�E��,�)X]���he�� �L��@%Q��۰�!�6���?�-Z�D�d����l��A�<�)-��ń֜؂��Ƽm�=l�f�PcR�>�Ӏ�����|R���qݩ�jc�Q�����������MM���Դ�L���̌lsV���K/y�v���b|���?��ҩ�vY��ζ8���a��P�c��E�v���X�t����0�[D�?AS��O�:H)��΀�N�"	H7�;[f�m���i`qK&2�|��"���6+�\s�^�;5�6���C�h��['�U�iW�6�\�?�Z�#
K�#��#�S��l��C�A�lN�� (۰)�W��m��Hj��G��m��n͐�ڍ�U�=~�2��'���7ՠ�M5����y޺]4ޮ�wB�)A�K�W���8���<�_n[S�$w���@�C !zR�B�8�$q���A�(ޫ"Ҧ��}}}��W��.y䣤VitbԪ|��n�*�"V��5F��8���KQ�}�C�t�j��rQ0D&?Ս,JlH�������ژS?Mj���gW=��v��3l�{���j�b=��Ԫ֭]����={_�~b�8\e/���k"�)�����sBY.�R4��_k!��Kq<d�k���DaȠbB��%ד�x�)v/��Hm�6̲����V�Kwȍ���(x��u���d7����i�����1���1;6>n�S�6;3k�z��k111�0?��>l�GGmbr��5yA��qB�� ��xt�+3��˗��c��@��Ј��_�����6Aюa�(�̰!N^y�_Ɣ��JQEML��U�l�M����'��Ɉ��T�3�������2���~���SE_�jnq�������X�8�*^�B�x�G�F� ��Д&|@��1NXhF:*�*�_�o�a�ݳ_��*U�r���A���k�р�#�j��?Dhw/4~{��za�PW���x��ibqZ�v7#G�#�#5^@����4��Im��O��W#�ڢ�ف-T�m@�uh^�ʱ��Y[���.���֫�=�-ݠ� �����^΂�ϝ����O�<֕��:QO�(��/��?�B�Ɗ1y��;����*qr^Y�P9G�ڼ(�~ϳ�i������ju�kR==ۨ�Q�Y���2T�O��ҏ@�=T���BgzOU�!�di:�tpp�T��kv��Q9�#��O\k^x�]q���Ï���)gű{c@S��z�Pmw�:��Hj%P̯�S����fzG�&L��8�r�E܅ʐ�����1�6f��(Rvt"/�j.>'�,@�ML�L�Q�	��ĸOB=�=6<<l�֭����ۆ�l���n�:O[�n��]�f횠Q>t�7���n�1vEG��C���4��
}f�D3:�'���w�b!�Y�a�'���19e��.2���I�3���?�ͤy���T���kj�p�]��3�Ew�'����on,�XE�d�֐g�Tm^���o���M�de^��J��������@�qY��̮����F�1��-�Ҫ&�QZ�zR�+B��1����5�ܵWsJ$V~�-o��������wۭGd*�[�����=�Q��ʭ[lq�fd��^T?"���۞s�v�iCV���j��L�����=����Kΰ�_�۾�m��m�n���Oڼ�#��PA��sw�S��egl�l�8 %k"�"�ع�^p�۲m�=p�mYS��t�]�s�]�k�]�k�]x�F{�郶g�ݵ��Z�����%�T�#�Fh>�YC�Lz(+@&%�<���P���m��crIP�:3u�*��}��wG�X��9M��|�P[{%ql��tt��{��_a��z�}�7[ud��l�n�Ã"m���h̬Vw�q�]������O}�S�L��8:�yZ[��K�4�A�C!�s=ֵ�VY�Te�U۴q��>s���GԦ��޻w�;v,��?)K�ZԠ:�;d��a8��� ���9��o[���J#5�$h�q���R�|�����4���#�2*.y�4�7�N���AnLj k�D%8���ƒ�uO�U@��W�7x!��א希]	!_'���W+�lhh�}�]��"���p��r�a�ۣ8��S�V�������m��C��T����9�z&�hJ�t����r@�H�e�[��{<�����6�v�$Ҳ�O��"�qx'J/�/P9ֽċ4'�)�-W8q~��1�o�'��bgo]c��d�.�~Qy�뙷������'�ٱ�f��ؔ]}���뵙���U��p�z{�������I�k��=Yn������=�����6���i��~�x�,H*�8���OV�W�
��qّ�Ƣ����{օ{d��ʯ��������g����K뚳͍�����|{�g��5���n���v�aW�g������lO�x�ݱo��z�!�̵;�0g7�7_�]�CO8Ӟx��dǈ]�uĞp�{�����gl����bf4K�F�6��ٯ>�)��i�7���v��6�Y-��˯��~�Y�ؙ�7ۗ�v�=~�N�ݗ<ўv�.{�y���n�'_�ݞr��h�N{�n�ɍ	��U)uQ�\�1�.�I+�9��@@��1|�t-�'�b~����(P��7�J�F�H�/�A���J��MXOc֝����|�w۶�����n�fS��m�q��>g��������s��MNN�Yg�e�_��'>�	_e.��G�;\���F<��r��H9�9�U������i��Ӷ^n��:Y���n�l;�:��ӫ���|w��nw�y���}��C�.-�ؑ�a����4$~�{E�	+��d�y�q��/W9�t�%�#.t����];��6����&�AX���i�4w�&�:�����R,��蔿� ����p�MLL��ĤOL�֮ӄ3d��������3�:�eٙ��U�Tc2b"�.����n9�C�==r����B�`LNM�k�k������:a)�";�Zksk���8��`�Y�NФ���f�
�ō�T&&&�^��ǜ����'�c�;�n��.�oR>bA9	�+�ң���?�|{�3a��~�}�+�����j���=6�ė�8*?�c/�x���3��'��ӎΌڝ�mN�ig4�X�+���_|�S�){v��z�<�	Jʈ�b�\6�		�`ٹ=�_@�}{��YE�̂���`�,���J�wf������K��fgh[O{��Ԋ|vޮ��|۠RM���L�c}ڮ=Z��?����w����U�l�D�]xҮ;8aL7�W�<��-���\{�P����q(�j�I>)������ �)2[��M~��h�6�O�j0�-T���-�mt�nG�٦�K5rr}�z�W�[���]Z/t׭�L�{��U�m��#��Wq��
�5 ��3� Ҕ�F�1�[a`��N�-��LVȾs�NМ;��u륟^^3bkz5}�=n��{,����ĵ>}�}~L22<b�i�S���9r!��8�5k�x:�Up(eހ.q(8PN��)�@�pFZ�������W2��/�0���)��q#_�+�Vk����x"���K�&#Q^\S�0������/�~�	'�苄�r9���?�>�Pm���&�oqJ�d8zJ�Y,���I.�H?�c5�mۺ�w֕*ߟ�<��?DNd.e~�grc�E�;��p��҃>������?�ð5�ZH��a3n/?N��)aIz`,5����M��Lm��ɏ=�񏶾���<;�K�am}ƞ|��֯]��cv��1?�������~�>��g�k�?����>�r;w=�Y�'[��.hA��>9]�r��= NY��'m[e�v���@U��$��uS?MИ����Y��(������]%p�=r䳽[�c߸�&e�}���=gj ��&'�U��ǜ�G�ü�v�A��dW�m��O>�J��R���Y{ǧo�׽�3��w|Z�){��}����w�15���엟�,ۆc�ލ�^5mǼ���sLڥ(���{횽�'������/����Zq��;�Ǖ�;�����Z�1=*Q]���?�L�o/��~�鏱uݓ�͊弐{Mre@e��'��t�2o����� 9�2p�'�V`�7#憮��N����ٽ��cUM�E�k���U��E&��j�s�e����������i�����0�"�������O���؏������O{:�`6l�W���?���?���}��>[�n����zM��~���5?��P<?A��E/H��{�����y���|���9� Af:�e"��d{~P�x��	a���y zU����1�C׊g�IƑ�T�¸��S�������e�z��nh�0?i#�;5�V-���e��L@�?07?�ΡÇ�>��lܸ�!ގ\@�r!�)�ιɾ���Z��ވS۵�e���s��A���r}��yzsu�JTw��S�`�֐��v\`��>E��z`�f�~���ۘ�+�8�v�_�r��9���=���Ê�ڇ>�9;V�^H}�O���a�ج/rqT�����Ox��ӆ���/~}���m���_z�x�=϶���3o���g�S�ڭt�WK	�7�����̌�W�tك���HM �J�J�4髇�lT��͚�.;{�j��,�I�ї��T�x�w\w�ʳ���Ǟ�]����j�������ۭ���١Ɇ�Y�/��������>w�-Tz��gm��=�|�ڬO ���G�3_B��I8��a��g�F5A~�	��}�>aA?:۰/�=m_�D�O}�jr��]ök�&{���=[�y��o�u9��>Q�CP�\�8�X9cPi��]�:0��$E�i:�x�C��@�'2d�`�(9�	#	x�gjE����.��y�l곑�~5B+�}5Fi$6���sα�����G?��~#y�S�컚���D�s��U�Bhv��a�^z�?B��z�_l�z�|�B^<���
{��oO|��F�Mqf��J���S�i�f۷o���+W��j@��bR�N��'�0l����1�Qm`_�x:����1,*h�EE��R��zH��� v>�5i�nv�-n8
I	�h����M�*c��-4	�-����������C �n��^�T�8��h~y�����ݼe��'������St~��vEӎ�1��5B����Y/�����5�2�;b'Β�I6�|D�`�x0_p����M��4�(�e �~��e�}�����z��6�I?����׽b�:�u{�S�EO���-�YOM6�z��w���+�Q���V�<�^u�i�܌�,jB��,����Y?��B�_����\gO<w�v�����n-�5�����!uR��mFx���~M[mlZ3�Y�A�̼f��ݯ����u��+��i����Ţ���?=�qڎ-�]�u��u7h���=�b톴Պ���M��̜^��j���������G�.;�lm�D����d򤳔�{����	�������
\M����S�A���Z��R�v>]��T�G��Q�cN��rE�@d2�pU +$/��q�C��H:;��G��`�QTz{�;�CǦm��2zg�
5!X{��z�w��o����o����/����G^�[�L&�{���Ϳ�f��_�{�{��2�z���7��ː��<Մ��/�a���������/N�c�mT�i ��A����V�[����#��AC_�g�T0�2_�<��%�.�+�gE�5�B��e�O)_J�x�� !S��2lA<�J6uqʁ�%��ܼ;c�q�F۲e�?<�r���.�u@����ںm�Ǚ<����Id�D@c�^u�n��v>*�ᑰ"��h[�)k�.�S~����݋�v�9;m�Ͻ��޶��ؾ�f����ﶉz�{�I�大��1�|��k)u�	M5u{�w?ͮ�5lCZ8U�(\��S����LtiѩE{u�aC�$Z��㻦mQ��~M�|/O9MHM���;~3<h"���`+��>O��H>V_���p�MK�3��ۥ���~���ܹѮ�2"~�/_���{%��Ԙ�K���-�uw�i�NqCJ�]3CL;(P3�4�5h7���΂��a���W�f�4@�(E���m�/��Ԡb������G؟����^�]v���in�����<����O�������-<3/��|+��PbXUGp:eg�4%�輣[�fBj$#2#�������q�@������Y;0:���+�䴹�_�����u?���S��TwH###��ip`���ӵ3��
۸q���� �p�v�y�G�v)��ˆ4���^����Gu��N�Nm�?�M��E,���e���S6̫wJ:�g�x�#W��𼈗WWд#�Z�p��t��ry#-��!ŋr�X����5�zB��������֭[mhx���u�ÇK���;>����p��m�Ɏy[z�;k����{@)�1�@8�=̶E�l�)���t�',7�M+P>� ,�TOw�h���ڍ��i��e���v��X�����k�"����7�e�a��'�����8�{x���m|~F��E���.�-=��4y�SJ�GS��#��/�T~�J��g?ֶ���7{�E��[_x���˞l/��|����K��ݢ��.M@|�\2���A�PE641Tyn�2h�v��6>Ր���}�Ŷv�a�ٽ�z+�v��e��eJξG���z[�qw��f��y�y���C��fK���F��M�XM�yo�ˆ4���f��k�*���g�B7�͘ )����S�����^u���vᖵV�lkF���Kε�`���M�k}5���	��}��@�ë�+��v3�7SD����I)�W9���-��h�%�τ133�;��r����3D{<�y����~����g>���������W?s�D�Q�Ӟ�4{�/��~��~�.������}�o�?�foy�[�{����<����?��=�\����?��I7w� �2�N�������Tq�1�5ہ�y{
�,7���ǡ	��D�Rd�G�U#���dڐ3�Q��� ?.@��(��NG���;Հ�u9���qT�{'���1��A�[�6��k `k׬��۶{��k�Û�Q)�D��x�����?�ү�����F@�/29��E>ub����@�3f�����2���|��A��u{���]���=�640l�ߵ^�Ђ�}���66)�7+��;v��'yqP�&���[�kn:h�C�v՞���l����j:��h�v��؋��b/�p�=�3�:8l��5�p�f{�������eO9�_��PY������`�-����D��ib��������/�?|�F�l�쑻6��.�`�?g���h����?��b��A;2[�yյ��-��=e���5���n���pM�8ok5��hQV�$V�ip��h�;/õ�P��;���/ϰ�y�(�Il��n�����i���ƽvˑ��\���Y�����n�g�r���(|(��`�|/���+3#V��Ke�N�ey�S����V�����a��ukl���nX<��Ug�e6J���G}�.�~��������}�������3�����߰_��_�?��?q�<X��ܪ�u�]g����k���۷���%��Ğ�������>��D�Lfʦ����|��V� Y�zs�=�O�y���'�*�4�����'e�ID]636�v�!�ASL8�/��_�+�O<c"�v/��ȱj�����+�;R�]��O3�^EsB��E�ɶm��A�x�Jh:� �4���)�J����ck�F���f���}W�\˥��Y��/�}���l����/��jv���>hG���P�L��$�u��X�4l�MȌ6�����g���j?|���ѧ��M	_����R��'g�_o;j�|�Q������ջ4�M�'o��_���Ǭ���b� ����gL���� E!�\�H��������=���g\��n�W�_�s���D'g��T�2m��w��5{��v�f����N}*�dj9{�߮<}�R�v�ظ���cױ�����<j�P�}6FN���"�0�,-w�v~v�����`?�_�7��c���o�VGg���i�������>j���;/�� ڰ��� �ma��J��ʇ$�%(��DLGq ��!}�<�ufQP��������c��O4_���|�s�������|��v���ǯ��}�_�3�<C�x��b���������������غuk�%/y����/�����k�s�?��$�j5�R�K��+��{,�.�� �@u,$�b��!�0l ��v�Ѝ�w�A�|�7+����6������Q>����j�!{	 YJ�
���:X�Ŏ�� 4�v�	��w �D��M��A:�5�:��B/� �l�j���54vT���Y�`K�^�2�@2���%mr��i�Y�#s{��nֆ�n����^��l�@�v;�w٬�d���I@���5]��;�L�OhƂ�hR?Z���������u��)��.���F��`!ݰo��~����_z���賶orT��?����]k?��O��}��'�\�=^�0U�_�͕�x��q��!Li�{�^W�E�o�u�6=�m���.��k7��9��S�O|����n��n?z�v޺���Oi�S���uUv��n��W<Ӷ�_c����/�`Sԭ�֖Q������>)�a��u7�Z�x���ڣe���O�a �ܒ�פ��Ԭi�V�ٹ�i��������)��f�TV��O��:��V\1� &@ٿt�:�FЁL 
��NYl�+��*�~�m6:<�Q<�z��)+�O��I�nCC��U�x�ccq�FL�'�ZT����v�g�|�GϽ ����!߷�q��w��7���-[6o��w��e�&�T���?����|�>������y����/~Q݌j���vt��dI��h��­���y��E ����H}N�l��ϢHs�~ؽg^���Io��T=���V�>P	�2�F$@��s��OlB�'���r߷ <]�&���"A�� .><ņ#f��]�Ǆ#���;�w`��@�& ^��n�c�b$���MxJҹ�w�;$��^���/_�+��X��u�p8=�)��6�(%�J ke���F߅M����]Kv�]���ӗn�N�����3{��d�7��ث�eo�H�I)��?��wOH�'Ш�VS����}^>��eC�I�4P�����U�Wm<e<����.���t�!?*?;�rs�u\��c����6�ߑ*5�j���P��=�B��Z}�v�hr����c���׵⊗�J�*�cv_8������U�j�uޙ�ۯ|������go�g�����"���{�=n�&c��ܦ-�}ru���i�ڼ��^��쉻��s�=���R���55\I�Ԭ2yҎY�W�x�1����1��d<R���u;6�cܤ�
��纂\�<@��>��1�I���&o�%���9�gg8���eٽ<tXq�َ+'a'�4�	������������/�ܾ�؍7�h�~̣�Moz���/����o�3v�a��ݹ�G�7��O)��l�&�O����&��z�_����v{�߼˿$H�w�����D�h�t�~�\� ��8���P;Hs��	F���q�&��1�k�-��+t�qER�t[��<1R��,�}{FY�˼�͜$��i��ʞ�8_�������d���~�}RF/�a	"�'�X:�&ot;���K�EP^����	��h�'�T�s;<V�/�q�|��i٥����hc򻼅��и�Zl/���9��B9�u���	]��6U��|�v���l�����vy~Q�U��Ŋ6%�;8�0���zI2���%}:�@�4���=Vh1�0�/�k�r�>���u��.{�_�}��v3�V4���7$������}�ޣjT�=u�&{�w=���G�i�z���-ϼԮܺ�W1���-��w;�̓}f��.���ءYۦ��q�����췞�h�5<isS����c��#����6���y�SR ;@���+��������~�ݿ8,�T��p������%Ω���/]�A���P�#s8��z�&���v=�+��<��Do��	;�����wڇ>�!ۻ���io}�[�������������~፿`�\s��F>��O��?�q�	qT��7��&���W�0�9�>�k?~������;��$�?
.@^&���b5KYv= _6�2�g��h�4�ڠ�f*�zI�i~�r@��p�zt��+�<�/���#m��|s�o�>���=,����o	Hm��u�P�c0��r����B [ɟSy�� �>�"�R����t]@�hG��1��%�;�A�Ȯ�b_��>���-J���_�Q>�_
S�qz哎&����5�f��b*'�����4�ǭ�����?��V�#��Ś<d�
Y�W3o{�'���^{���o���n�<Г|n��
�ą�}q-�K��,�A0ԨHX	��ˑ"�o�O�=f7�.��59|��;�q���=�b2ewf��{��|���Ǿh_��q�FU���q��h�;8a���o؛>�e�{�bI~�������h�����Nh�y�����kn���=6/G�m5U�����q��v5��k�V1�f4��Z��CvW�V��U1�]���(�;��&"BGJK������"�Wa��'���cD�w���"�N�������g�Io�{�A'�U;���������۟����>�9O����w�	񶿰��_��qWn��������y���fw�s�O�`�f@�=0Q�Ӈ��_��t��d_�BC�v�����(��9H����cn�A������0HW��[�K��R��s�(Z���r�?H�O4��
��B�Ss�r��:Vu-��νЭ[��L-�/�� oQ�v��}�.N 2��a��x�}��}�T���~�Z@f��2�$ov��U����(;������E
>&�^��1��ʿ�J��E�D���+w�N�MS��o_�ۦ�|s{���s�����z�#�ro�e�m����ql�����ƀ�v���m�:`����m���yd���p�����ݠ�9[�#��v�k�Mj!O��:� ׍�H:�d�p�И_|�m����2h�AO�p�Q��DJ�hkװ�ڮm����19��v�Myu(U��	5�;e#j�i}����Ƕ���f���v���Z�i�>5�Z׎i@3��I�2�]CU۳��6k{}df�<v�8R�c]C�S[�.iESuW�b��U���z��u9q�>�(̍C��NmQ�b��<�#�:�_i�W.��x��&~�SW�*QN�����*fe,��h�M
Z]N�-�:~�E�u�ӥ	���ٲm��Y��~�g�`_��N�}l¶�_g��_����g~��~v��a{ғ�d����g���nw�uW�H�:纘���t��bŭO|����_,����f�s�6�[��lЊ��6n�e�ͫl��;l���v�-w���_O�%.��6�������?~����+(��@��P��%�G��7D���}�*	E�Fy�x6�9
Տ����ٳP�������_���z���W�'�V����2�}�DL��I����b9�,Ϸ"d[(����lM_-p
�O5�rRv�|�ȶ�}�.����FT�zk�vh���q�5���,���-Dr�M���D�~G�"�p~�_��S&e���s{
�i����u}V�?���S�6�M��z���J���Z�͢���1X���6-:O�Y���.�t����f��t�2g�x������E��_ǎ��H��ap�G��
�>��ů6�ыo�|�Y����PB�(e%Ϥ�Gr�=�w�Kίn�Mv۔&����̬�5Bq���yME�L��0W���k��L�n�o���}��	5F��D7������pu5I�A5m��w�r�>zׄ�tH�pM|�9��Rk�~���Mf7[�����ݏ�������W��)Ѷ�r%)�O⩼1��tـ"�j1*�<��>r����g����j��Шլ��U�������O�̀]Xy�I<�{�|M��v$P;��"��xz;m)�(	���V��5ڢz�����%�ᅀ���Li~�"�t��Ҥ�ּ�ET�:�Zb��	hv�EY�9e@�Bv�L<8Y&訧��7;@B�F�9��>�zW�&�;0w��2��Q�O�q."���]�pP��$�.�+����#�$I6�����������NRH�7��w�/�6:S�,�Z1^�|����s��@���r��97�g�鲻���m���OvD������8p��)u3���N��'�0^�o�8M����EV�.���{�!1�hx� B~1���-��ݫ�n�_{�w��~����"��z���A�fIvɺ*U��)�T)^��݊2�����Р	�����)y:��#��${9�R*q'�&������'�2�v;&VQ���!�͞�����T�|X[];�?{�_����3��O\c���k���^g#1)�2*���lp�������t�����R^�/�:�#��n����{��{�{�پ�/څ>Ҧ�#޷w���	"t��7WG������J͠�q��8�W����A1���Æ@t�S�i�n���X��޺(^̦=m9��xt�0��|y���9ye,AG^߂�v�;�$@-�E��s��=C����v;<	Țsw��p��q�5�7�XG� WamG���E�b��,�b�c�]��wN�/��]s�]����Ly�JP�'ݺY���
Oѩ����L�X�%��?���:��x�O!2�U�H$�,�Xh��O[]g���Wg(��@tsp�PR�)2�1Xs��H���xVNЁ��
9��+e�n0JSb���ǡ茢	'�����k�T��Oer_d��;�b�@i1�dpDlȃ�y�}���n��~�Sv��?i_���N]�j�ң	z������/�%О��)�S����̴����wǭ���Ƨkv�]����x�%�J��F4/��xb)D��� � ��M�"�H�?�[���Yѝ�Cj�[���Co�:h�Z>YVan#��5-v�|�����@S���u��͗��������>��p\ɾ�,��:GW�Z�����������q�i�d��U*�⯄9���Y"���c�	3fȴ��wr��k�&7�3�ᅀ��t�����o��Tb�2�v���Ӌ��gZ)h��|��K��w[Z�o�P.�����;��m��q�^��N9~�kANX*��O@�����8��еJ�cc��7�/�ӯ�HM�V7L2N��#&e̯��f�;��2(�/xD�ꏾ�����<x����_��n���#�"A/�hF�I�y����@�1y�6!�b"vz�I:�.a"o�D��-E�/�֔l��� ~���Nc�� :��q'���-�6m*t�� 󉱌N�=�_�������}�e�Z�˽ԩ�p�B��*��8��|�kZ�xITf����r�1h�� ��B��͋ix3�f�⑪ t��~���mŔ��Bk-�	�
��<�I��T�>Ƒe2�ڿ��x�y�A�������Nv�o�uE��BQR��ݕ�Bh=PDZ��Y�c:C�c����ݐ�(��յ�/��Sx<eh�lD7/�S��}�}1�N�
{xlR2��Lo]���h�zc:����;%���0���';��O(��I璳������&�cG���}������a�ڧ S�~���[��ӌt��9f���ǵhZK���$���`�%$�y� �ɇ��� ���An!/v�	@�ΗIf����8!���`��~x6__৺����*�fF�.���V���R!6�S���y|$KX��B~�������®�.F	�<�#i]K���:}�[Ԥtl�9�J�IK��m���kD����� eA$� �]��u_Y�́��#�v�M,���rvm�༱��O]�	R�_'�#O�<:?����K��mHiR�n��^.Ѵc��	��9o��Q�<m~dUU��f_���\i~zb��qet��w�T�t��eԵR�M-�s�G�qi 1�d:&����[ň�<_�ɲ~�ū6�Q>�0��9^LH	���e�v�'��ҷ#��r����C�U�_�~p���n�ƾ���Ҁ���Ը�:� ��B�H7~<���f��y�G�*��I2����]����?�*��X֛�C�T- �v�H>���QL���J@��j��W������ن�����Mr���\�'"c�]ƕd?a�Yb���x;��o���gtl���4O���4'��Yo|�d�73L�\�Z��4��wk�[�&~`�|�~4������-ȗ�t#;�Ub��xO����8-�6QVnE�@Yx�o�5��(c��۸k6�o����i�=��n��~�����kL�֙Y9g�@*����!:y@9�29�\7��+8(�Pp�sp�(.�R}9Ub,/����E,����~���[�Vá(ȝ�����@y �Ľ�<B��]���������K΍4�g��ں��h%�����i����k�6���"?U��|���3?�S6>>�7��Q��������[v��wP��6�ՄB^$KbY�'�i99�x��(2����L6=�l��D��%wL�a�n���P�&[P�	y�ǰ��jӽ����X9I�P#r���]�2����w���膸#t��t�t�o��T���F�*�ݘ���Q�ј���h1��q�~S�r�N@���/~ho����s�vYR����4ǫ��vJ'��ܧ������ 
�����[dm ��ثyd�N��z��ޡ�D���-�
}�$˥���ס<}Hs9.tWe���Pm��ؕ��x��Qa�$���γ	����qr�ݹ}�䠔���#SHy��$. �`���w?+��ج&6=�~;8����1k��'�3.�ݜ|~�S[��}j�Λ�k��6S�7��*��V� (˅��2�dj|g኏�w�'�F�W�D���=���>����o��<î�����7%pYV!G�vf�^iϡG���M�	phr4]��UkGm��_Μ��D��OzDϗ�Z�h�Ѩ5lb옭];��Z��SP<MƷ���O��t�O���؛+uEp�.�BU�Y�%4� 	�����DhЭ2��'p����MU+x�84$G���wHvy����F8���hG�X�g��2�G���6�b�B�5�
A9(B^3��Aay��Zw;���ɏ|m��ɧOQ��Gr����|r��p���C6nԎQ�?n�o�6���ߨ��d�3v��§wyyHn��&p\N��0�l�i��/��u���2`���84M;���|�)]����öyr���f�Fi��)��'�.!x�&!����I	��VQ� b�%&0���o�N�'�d(�v'H��O���j��ԋq4b{��a�6kGT�������ޜ|^�i{߫��]8~�.�V��kteL>KA���P��Ѕ���6�rut�">��;	X��y�u,,٭#�����6�+9f2ڊz{V!�K�*&�y��>Q�EuH�ܤ��j����bc|���qr��R�δ���G�|�`������'7��0�YL>	�
�0A8(�-]x�����r�Ί��4*r�wy���q��lG���)�A��l��G�\ie��$ʓr��ϯ��=!�#�t���c�\��O>�YJP9���GmS}Lch.v>"��}U�O�ϳo�>;k�Y.���W[�?�^���v��5NxS�7jt�$:AYnn6л��m�eS[/�%��OIUݦ���}�����b�W�n�oۏ���2;�(�>6U�
���ʉ��īd���?�O�5��y�:�F�+����c��6v>����ƺ��{��kG��YU��O^�$M>����i���ٺ�C���m�Мv>}5�G��#N�M�t�r{C .�D�x�d�'%;���l�L��<Q�c�n\��oZ�����޾�6͊�g�Ն�3R��V���+O>M��N��R�(��G�8�L�.8�Cd�kr!疟����򜘹�ū>�м�?V?��2L�p�����# ���'%�еۀ��y:��N�?�30|`��'�I�kG���\�+����?Vm��7廬j_@�kN^>A$=�D����P�t$����	X��9���͵#���G��~c�\�;�ɇ�I@~?I���� .oч�� o��׎�:��/��m���,���xYlގ~l�N;��-X�5a�&�͓I�R�����V�#��1x�S�Z���Ʃ�aj�hS/��!�t!>���ڔ���mY�L8Q+��'>n�u�`�g�CL|\~ѡS���y�>y(��4mH����W����F�{��6Y]�/ ��/}��E-�fa���1�:��'38b�&T	%d`�⎞��������|㶯ޭ��ɮ�z�i��u�
g�Mt;*�Qn)��SFZ��Q���%�jpā�Q8�����6ȝ�)�kj��@:��AB����A�G�!7�o~��w���P�vn�����+3�*��A��{ħ��z���U{u��7�^�Uu�t�&�@��H\AE�V@䐌\w��xK�,����uU+K�kw�5�]��_ȯ&.��#��ڲ��V��MdWm��N�z�Y`k\g�n y �ZO�.&���M�ăOL�e/%�NK|�͓�V�3�����;����ڒV������}2����?��,#]�@a�����|2}��I�9���(�?���p�?蕽�ܣ�Yo��5�t�ڌ�t~�wYB���e��*�x�ض#m՘-P>#a���ˊ��ȓx�;N��O\��E����j�ڞ���)9_��ȹH��5��it�
q�E9�.*}��0�E��GZL\K��!I�!?w0/M����ˉj'���7��(�+Ҁ��� g�ϱS�o)T�y�Ji� 5)��ʨU�ℤW�WM�����p�
�|�����ĠN�w+/�z�r�B����O �t�+i2ӄ�O��mgf&1%�L��A���� �RF:�&�t���.&PB&�h��N�Zi����:c9M�&r]���@Yt5f�n)vL��!�}�~wGy o���Q�"�<�
��0"�sD���1�	l�����o#@~�%D�����7���Gz�)A�1r�3���˾N:�q\�8t�k�/� �Z_�#7�6�u;يҖ,L�@}�s�c����Wiht�I��%�x1�����,�F��[V����������Ф?�FȻ%�$��6)9d�����$����ědw�� 99��r�Њ~�%��%��	�_�*�w�U��ȝ�;P�E�B�k~L	���>:�+�m��Ծ�#�H����h�	��'��,�+�xP%��	d�B]k�Ȅ��s]Q�9;c�tG�	�4�;a��&���O��s�<2�C�`
���D��י.�f�-&�&2�D�dM�Y�#?����Z}TS�9��R.}b�\!q�#�@�u���uB��ײ@1��2�E >8ƈ��e���#��˞�B^g"��t(&����",�2�5���#�n�z*��n��ޟަH�f�{����=�ss���u�%3��+lW���=zY�11�����߈�H�T�k8����Ӟ	tH�q0���t |[F� �(A�D�9�1�F�(��wt�D�<Y�v,�f"�s-�J(��1�"y[h�l?�?F��%ƞ�"�ۏ���k��=�ڿ����m]��]q�N�]�ˬ��Պuʋ��Si��@l� �C�L���][@���SH�	��ײ����G��r%��8D:Pp;,n�1���إ���x��Na�Y���Pn'&�+��D<~�����Uz�zۅ.�_�)��KI9�Xy� ����������F�O�Iu��£����>I�0J��xo�T��J��Q��8!��* bZ�E��uM�2�s���G�*�k�@����Y��1y嵂�>��Z�v�Յ�v�����e�z�e����W�Pv�F��\}ͦ
��0tς�j�����v��m}}����O�2��)���Xr^��ݧ��:�~N�������������t�������@���X*Ħ��%��#}�!�aгȮi�Ǣ|���9�_�G����� l(�S�B�_Uu�=�?_ ���;�`�9oS��mp�%}�n��y���.�"n�0>����]g�tO�����*���5DQs[0K�a��"R �����e�?�U)����F��4����@x�{�Pв뉬W
��H��H����(���!]OL��7��:��T����B��i��(T�y��N�A�����wE�qp���1��&ԮG�	�p�vU�Z�Y�)�='�y����޾S��+��gq���Y1�SV�ᐏݖL<�Aj�G:�7;�Ѝt�a����@�-4�ߎ[�A��ŗ��m�߾���MsӶy��֬鷾�>��
G����Cﳞ���c���և^]�5#k��M��<3>L ����8H�%(�}����2��/3]����Q����?�}轌��O?y���>�f��_3�Δ/�c�����+�܎�s��vP9x�2�"�up|=,��X��B��O(y9/?@884�:���}������P�U�����z�Atzq��,���_��Ea����1K�E#]��b�E�W܁���U�r�Z��g�u�=�IO�g?����W��^����O��O���<ۺe���o���`_�wg�ơ��p����%d���R�����Cm:;�jᗱ 7v��TJ�-���q"g>������1�zg'�i!gr���	E+��gB�O�.� ��������hIS7�W��㠠�}"��"�eF�~�"1h��t�
�*�_�X�lΏ�; �&l�3��u:苜�A�Ve�C�iM>�l��k�\a|8�T�J�ՠR��Ś��Uz��Z	N`,�cS����n]+����~c�z�ě��WB�G;x�&
�@Mݶn�-�t�|��x(�~p�W.2c�ԩ��rX�?�M�(y(�6Q:?4D���+�~@�쳖kg��X�h��[d��E�"���<O��?����+^�2{�w_mO}ړ�̳v�$oEɈ��VEtUFt��՛.c`�\���@�Fߐ2vY��~�W����C�ݭ,���)�>;&E�VMe�E�CO��@��fJQ/t����_�m߶�������_`�}�]v�ev�g+}�m߾�.��B{�cg333�ߚ��O(*���.ꥡ).@n*Z�4����c=�~?+�a 	�-�] df�sUq�r�Rs���Ԍ��Uď�R*��L�#�&�`�z�ㄔO��Oq�n�J��[ҹ����чr�+Y��{�A�&�^^t���t|��x)t����_Fb���e"A�-ǁ#�0�fn��4.N�ޝ}����b�ki��[c��77�4�3�v�y���]���o��8?�����x�V��zJ��(���	B���odd��f��m~/�ɇ_���IW�
N��f���Mc��wt�����I|�Sѯ�E@��֬�C�l[6o�W���5�F#��Dy�S6�� }E�)A���pOrD�z��t��]�����.����[���7�|W��qE;�]I0Ǝ�����	��@q֌qz�h#sS6<7!�[Od�z�;P��8��2t��@?���'=����^k�_~��v�i�s�N�}�.��߳([�'�''�ԏ3�G�2Z��7<����!����R�8ݑ��V��Ȏ�u��g�:��zm��7�k?���X]��P�ˎ�%�9�,p�tR�׊�����1��?Ͼy�&���u��g�y�=⑗��u���.�mj,�\Im*��lff�>��O����^���Ǒ
��A�kf[�Gq�OCQ��<�[PO/hp��t�u�m���P�/SBf�N _�GR��F�^)�xK�d+�x�0�˭0�	�k_ͅ^
g����t~�溈{ ��x��Q���|�/�W�����E�3��8"t2/�@:�����F@^&P&�R2�����ϵf)�d/�IKՓWO+ʸ�i�Z�%AЗ�򡍢��m��.�[��ͳGl}m�����}�=�������{�ƿx��S��1}阜����s��6>q��M���	HL��	թ8;��>�v�UW��7׭]���>h�_w��ڧ�;���z��������/�؞y�3��s�vg�������/~���_�E���bD�.����s��l���W؎;lp`���Ɉ�}�:���?k��~{*�O��N�e&&�l��ͪs��$��#�C���к�n�7��m��^e䷐͋��	�9N��lű{.S�<J]��]1_2�6�W�^AO������p�Tz���lfp`�^�җ�S��d�����0쎟lٻw��r˭6zt�n��:����8JX��/��N�Dˢ�vp�k�_2�[w�e�}[���������k����f�|���{�1_��>sT����1�.9����M��
���RB��	��j��uv�W��|��W�N@�1תT���N?�4;vl����h_�4���e��L��G�9ڳ��zF$�R��(�]8`畔�ӄ������;��/O8������Ԯ���DW9ң�{#	��M��/��\�+��˞�=IE�Η�λ0���qi(iy��
/h�t��;�����\~6.\׫���h��������<E=.����:����Z�OQ׷����r\�ޔ1�0e�9]w��瞣��.��	�@g�aa$#^�t��~�����ȡ�r��fd8�Pw�_����'�Y���������/�U//���;��[�څ^hW\q��w�}�ho���E+�g<������.y�%����!^�4���߻O�m_��W|��<�ʂ������b�}��l׮��/��׈mݲ�.����G=����o>���*��L'�ɈL7�t�MLNjſ#���3:԰G^p�u�ǯ��f�y�]�Cq�`K�D<�8��n"������t���ynZ��	��i����6���a�����O��P�����!c�+>����M����I}{��Q� ?�(��I!����6'�d�p��N�m��������n�|���M�A$Q�jAڕ�4VL]t�������e�H��1x�
0�N��D!y�Ƞ$8;�*���2(���+�Ц��������z�j�栋)(�`")�+Ġ3/��=YX�#�A��~��'��Y����Y�d����]�r�U�;��?��߿o�?U��7���V�ay@��㏗�>��O���>����Rq��v��i��K����@�e�
l�Y�z���Mo�	ȓ�����y饗����e���)^���j���hE���'�r�Y{�'~�'�}�/\�C��d��L��֎�뮻�f��|d�X�t�^"S�<Q�tN��r �jņ��4�<�w��;��nQ�/D.8��Q?� �ӉU���_�7�k��a�+y!B�d0����r��n�b۵��Wn�J�JQ�9W���|'�R��(���?
a ��u�аBU�I�Vq��v�P��@'�k��s!d��j[�*mꕕ���?�2�s�A�tV,�SI�-P�^>��i�@��X篌eY�ׂ���D�\f"
�,q��%J����~�C �A�VY�uE��;p`���jE�Q�jE��"
-�˝`S�{������Ȋ�ess�Aա� ���?O������7m�d/y�K�z֊�uy�$���bJ��0��g<Ӯ��ʰi���)Oy�;���U)�4�_�/�;���1��!�	�I�N`!>L@#�qt��v�-���+Y��Ҋ�������$Q�X�0@��#�D�r��꭫]�_~������}*�_��٣F��~?�z)�a�	�R��S��Sbs�a{!G�KB9&#(c��	Eg����vj���x��֫��j���:<�0d�a�a6��ޕ��%�Vk�D��6j����P��i����-0 �c*�gNo�edL���l�~����!2����IL�"��N372����/-���������\\;_�����|�t\��U�f���ȅ�1I�O2�b���V{x#�Z��X+x�(#�9&bo?������Vu��O���j�>�Y�������c�����.2��A�D:���Ӟ�4o'��O��.��7����e/����/|��N�ArBw��W��@��=���e�j7r�ߗ��I�}�}��������/�?��?��Gh�t�2춾�{���i�'�����^��^���8�����M{�K_f?����N�_���.ע����T��;���䠻+U&�^�Α#G��{亮D &�	K�h�"�B�5K�c�m) lye(ڐ�d�	��eNX�9E�����Q��j��yӦ;��a |�ʘ�h_�ox:��v��qA�b
�S�� ~kְ����|Sx����|6�!cHvRҩ�b6Vi�}���;����?�������i�jW�I<�#d`�iR���T�ˣTS~�W��O�R��7�п��3�Z(�ܚ�k7���6��J迼�d)y1rZvvޔ�a�qǐ�	�Ii�
\��t}d���^0����y��Y�B�k���'�t]���E�<&��*ACR��" �Ϯ���Sg�u�mٺ����̴����}�ӟ�ɩI����~��[o��b�3w�<L���>�* �ӨQ��o�jo�����y�����w���	�v�y�_�<�p�駧������mn��Gm�ؘ�yǝ���{�}�K_R��h���V�9�~�O\'�'K@�R7:&�phx�����#�;�V�C��	�K@B)�9>�P:�H������\�|�����i�w��� ���P%���_�]	
�jK�����������U�O>�(�
\=4�.�O����Xs�΋�Ua$a�'R2&��Ln8�������s�j�֞ �X��0:49$�MI�Î@���4.L>�k:�2Y;d��.����	�יK��,�LA��ܒL�uJ��O(Җ��N�8.s��dP��%�s��������u��p�k�U���8����N)�_��}��_v�皉�����i���G��nx2����/�599i����I9U��}�s�܉�kqbJtgxх9o_���}�믿��f=~l�>v��|g�i��9{�m�~����Jd9���(�N~k�!U.����V�?�Y7`�4
������NR}��.p���V�,g�v���CW>=���P�$��t� 1�7 ��O!���oO[��l�P���Y0]r�\b@5��q}���!TإU�?��Qm���&9ŕ�P�~��`31��H��qp~�9�z8x\犂.wɐ�1��H�Yh�4�;ZB�-f�"?���!m�r�[m��Q�?pG�������
'��.�p��LnK�w�xd�?�3��"])���>��D�A\K&�ˮ.�I�ަ�;�����W�Y���%@Y�#�H������I�Y=GjB���RK_5*gN����8����Ǡ�?�O�1i��.@�:�=�؅�6m�m(��P%O��(4�v�Z2���'���
\X��j���F~� �N_��a"��9����܏�����	�vAЮ�r�g���#~�p@�����97��k�Z��୿��R]{E�Km���vt�)J�?�n��OB������(����� 9@�X�w����g(�%t�g�\��l�'p��>˃�d��e[k6�I�ߠ	'�2��$��Q�:�-h-��f�&��]���'ڄ�������|� #ץ�����@�՝S����tRN_����/�>�h[�K�?��EF��*r�m-��t���e>�!A`�W
s �nG�#��J�+�O@����NE�㛑seh�(��೤1' ���~�Moz����o��|�#!^V��z.�<�p��:p`j�٤&�_}˯��p�[��V��
]"�x�w�y��ڠ62a��q+�>���@{���"ٓ� ���L>YF�6��P�<T�:e����9��=�й��ŏ�H]^�R1W��9��{�q��)�d�z����HN��?�_�;V|���ı����Se�'�TU�M=���;�Y٧��u����G������RH�t0�8O)��s���Գ҇����đ�fG�W����� �K��b/�e'�v�~s���U�(A�8u�N����k^�����eX_��9\�7�h�����,����V��݊��uR\n'Xb�|�/� #1ʣ��nvZ��U�u����s�˰X5Պ���n�;����������_��������w�y��r�-���Z�y
���?y��X��	��c4�ɇ2P�;Ʋ�����S�vl<V���W1��)��$�y�G`�Z���PC~�g�/�¬K�lK�j&䘇���`����~��m)@ہv]s�5>��c�ܧ+:;vL���p_M(��m�����|��*q��硓v�#G2���̴�}�}vXIò"VR�;";߸���4�o��*��q�c�=�0���8Bwz�+$���/�4ʕ��F�(��@������V7����l;&Y�NgG�:Zu�&zĎ}�Ph�TAێ���\��������v�w,r���b���?�/鱾X�&�H�O��-0�pY����E����˯vq��@���h���Wd 6@ɿԑ���I���7m�@����$>��k �,B�ν��8�"4�YV"Iy~|�xv��(��+m^��W[_� x� $?;jxp��h� �Z��:��`��>���˗�� �*k0�(�8!�q��Ʒ��$Y�㴐�xns��������������|ʒ\���q/P������q�d;B�!ۙ�M�(3:)��~��׿{��wy@F6�GG�{	�Ec�-W6�c�A�?]��9A�Bh��I ����!��}{��7��W�_ڧ;]S� �����}������̬��/m�O Ш�vT�BP�Ets�F:^�s:���G�ZwHA���aj5�����.��)�W.�p_)��P�'M(�_�$t.��s�I�L:	$��Y	 u����@�	$�z�W���JG����]�Śt$0	��r:Hࢊ���6b/ /��.� 3�J�_�Խ�+]�)�WE+
q�
�̡K&�����T�׭��T�	K-C�ɩ�?���W���Hm8C��1,:�wI��:A�8��F�:�~���f�F]N��8 ���e>�l!s�<��#?�#�����o�Ѿ��/��>�����@f~Y��<7A��97;�h%��"+er���4��:��,tc����C�����~ {�D��lQ���G�#r\�}�I$�h�?�;�n�J��ϗo��;�;��ѯ��e0�rZ3�5�;���$X��RQQ��mf�ox�sϽn����)A�~��a�����%�須�r��W�~W�O�K�lO`aH9-.�̴"�H� �t�c��U5�kgw���i�Ċ�#�xJ*'��aPh�����*�!x��$Ó#A6/C�������!�IJ���#��� �u���a�kbN#3 .ɣ<��m�k�k~ĭK�욳��y������Q��"ޓ�o�G��9&�d����-P��/C9�,�����z*ঠK�ȴ�*~�̊�ʝ(����K���Ȍ����o\o��G���x~�2�=/��7����s�&	&
VΣ����ۏ{:��:�6���ө?�L ����^[dIZk�u<�K��<�V�.&�&�xUL�W�n�qU@�u��t�[�cpB��@Ww�y����+{�����iʞC�1~:�B����GKu}���_��\:���,A�f:�����O}�>z�5�h�����8!����\s͵������}]
��Ph����'W�R|'�@r&:C�3!H�k���i{\�+m���X)>00lk�n����64�]�������q��ln���-j?Gj��4����Á����l��n����D�ń�,B��������$���e�9_�L��Y�GE��\���� �q�)����(���P���鞦z����$�A���nF������N��B#�.�&�+��T���l@���c�#gY����3r��{����g� ��n��� ����H����s��MBՂ�h��)dzp�L:����bA��7/��$��EQ^PL�m�Z@��	f��$���^z���o���K�Gq<���?�?���簀�>������_������k�_.�2�|��i/�L�N<��k*�>�.#���P��b�Jb��;b�JBf�<O�&�S���lM���sѓ��@����n��ׯ����S~�Z;2:O�z;�
���O�s���}�3��/ߺ��{c׹\�!G��	�Y������n>t��麻EW��Ƽ�;�jR8g�{�X�ro�tAS��
�!��2��+�8h�]�)����~�����n�][�k�/�����/����&�f'{�2�u��2�(M��a-,Vm�g�ƫ�r> �Z*f��O �"��ǃӱKm�N?�\9�V��b}�������x��z��ip����5v��g�ءC�Pc"��H��;�p�n�1��^��O~�,�M�e��\N2�>^(���RJVz���b�8�M1��'���	����Ǔ[�������i[
*Kq,��:so�Rxۑ[}�')IGL�8�5C��̳�`���[��34��J��:M��i
�9M�.۶������0~�u���+�P?�ہLȐ�Oe��4����`}����mؼ��=�<�������)�QfV�q�Y{��z͏��nΰ���!{�2L4��v�?��}[|{���w���0 �'�'���}ex���^���r���G�����hzr,���&|Q�G���ӟ���w�}Q���������%�����yí���u8�L��|��8��|��F�mߩ1]�m�y�ۄ�/��*Cv��7�|7�ދz�T�Hm��v)���O*�s�Pm�Ff'���u�A'~A��-�(a����z��O�3��O 3�\�	����6����yv�؀W��3x{�Җn�a5݋�vx��w��<fO��t�`�z��leˠ�1����R?��eH"���zٖ�z�}��O����5�K���kc`����P�Y_�_�6!u�{*�mA����:��x�%��+��e��[S���>_�ѱ�ML�M�,��l�&�vlz�ƅ��s65[λ#iԻ�6��3�V������-��Hs�ϐA�e�<�"�����o��Q��[A@�	��)�d!Y҄$���N���d�N��u�+ڂ�D�J�;K&N&yO�F�<zjV�c8,vA59��G���Y����X}�&g��6�0mS36՘�q��+u��̌-ԅ�A=.�d�:tm�>�gi��=Ɉ]��@��!��"�V�D���AWJ����m�qRԙ�'t��h"�,��i^N|O�u���/��������O}�>�яo�4������6d���W��~���ēH<`���n��{���<��dƛx��CTa;v�T^<���:֮[�oY �^<��.�m���K/<��%�{�����D^������>��Wuq�\�z���.=hR�#p\�D3��@p�ˏ�4�g>�_l���w���7{8/�E��\VڃN�kI�n~]��(��1:P�m�RI�n�RTeB�+��un|����1�0��X��A �2�d�(�Ʀ�ɉ�l�t�0�q*����;!�Z�AGD�K��%t��(՛U��VB��
�Y�J���*�.M<]ssf����3�ib�]r�@_���(���-P�\�)9� �4��h�N�:V�;`x
�p@]���	�
�|��b�*c����;�Hp��2r���:nh����Pq�<��ڬd��*j^�kA=!�<���B߱����EU�Ϣͪ�����i�^�?�{a��C�/�!iIn��~s����:�Jy1Q$T� �招H�K��e(t;���:���CA�m~\�3PT��3�ڹ�~���.�袂�����������ˏ�|�S摀����ۭ_��W��h�\{���a_��W[�jSv3,�x�!�q���)p������~vG��.7�y�o �v
�F�tP� �%�_��8m�@�8���5�W�=?ez��C����v��(���C�K�%�T�ʒx����1rNЇ�8a֏t�/����]jO�"��r�ZU�1f��~�JpB��/eDX��-X����_�y�##�|���m�H��T�%MF�1;��$��|"C���� �E2�tᔘ82�1����>�pQ����9��X�,���Gu�Hյ��t�F��*9*5ݜ�҄�.9G9�n��P�&E�8�pܮ!<���.��#�#��#Ð-t�}�l�s�T���JC������/#TJ*4AuF�����t�G��	lʟ	��&��Ё�uBUT��B��E�Gv�y|��qF^j���:��_׎��Uߓ�%G��yB��5�m�-�'l?`p}��Z�$}�k]2����α!��.��i\��l�����v�=�{���"M<�N�ǟ��.��?�};66�|��L��Oy�S�Ϛ�5��Mr"����G���k��oY� r�����<]�_��x��vU�K��cG*�����9M���>�7�����v��x�7�y�&���%6Ar�a��]C]v��ʵ7��f���h�Ʃ_麍Q��J���8t��� �Բ;A^�]���>1�W�˕�����Aa�g��8r8;BC��R�I��9�>>A�9�q�N"h�Ф<:��̃r�Yɑ��� �r 6��6�U�^Mqn���@��$k����G�{�Q�J�e�.9�-
�n��^ ���� ��x��BO\{�6<� L�/8��Q�ip�� �Ӷ��y�O�>������^�+���ꚰ��/�S{�x
UGM�9뭫�.��>�W޼�愄��U��KX���j/�<���g ���[�t']7����Q�)���(�/�<��uNL: �=�a�O,R��P��d�Z���ŽBw�.b�$ĕX�+'��ۤk���9oㆍ��7�ў��';�8do��}�Doʓ��P2�7������q ����>�ۿ�[m�㧸+U���:���K_��T�a&>~����.�B��O�3�<˞��'I\V����n��E�����R\�);�N��[��������y( ��sr�-h@)���� ��џ����x*�-�</�5qi���?��y���P��ړmE��C�܆��
]����|�^������l���=�����f����5��V��(�|�UVJԛ*a@� %;m�����B���lOs�a�pB��uDY��s�r�&�>�sp�=ؿ�*rhچ�l8wB���f��G!�">{ν��*ۭ��q�L8��V}ӆ�69>��ӌV�?J�]���?U���+DO\+t�W~�h�$�E:�����h��&�6VY����˔�!i��H'>I+��v�NB�*o�cD������)�I(,����Ӽ��~�p����~T}*��xU��>?m�:�Nﳯ���_�^�{vʏ'ei�����C�.^e;ζ�L�֪z%���Q[S��mö���׽�>��P5��a%蓢���}�T]�*����h��T����?��Kw�S;������'>�>)x�����r�$�ń@�P���_��_�����/���Q]&vI���	��H���f>�7�?��O�-7�"6}V����푏z���H�m���7�S���mټծ����u�ɣJ5v�.?`Gȇ-Po;�uV���k�� }��&?����sT�6��T�]���/~��J�_��w�X�|!?��Q5�fq���i��Z���/@W�b�2�l�8`[F�~n8E��$SD�Y^��r�Zy4��f]��/ʫ����,�|y�3�.N�Sk��δzu��a��eO�\x�Tۘ_���צ�g���=r����&�5RVtܲc)�S��m8ң����~�i�B��9��A�TD�ovx�Q��:�EЁL��6��kp�=пY�@L�/��S�q>"�H<V����4��Z%&�J��*I��Á��'��K S]������e�J� W�2�tVQ��䧱ڡ���b��:Ї<���2!E�G�A�S��z�MRϋ��u"��Z����-��1�,.b��63ϊ�>bh���[z^�nخ��{j�&�w��ӥ]#O���T!� �����<J�����0��
`��4?jkG�����m;��^��4��I:&l}����?`��+�����Ҧ��S��P�2��r���o�i{�^P<���'	�#������{���N���������c�&T�'#��4����?�3���*�=�\��?�}��m ~�W�p)ї"�������xY�J��4>q�\0����>�=55�G��_x�t��]K�Q�e/z��m�j��v&�uJ)O>!�/r��4YH;����ak<�6/�Uu�yR�Ϙ&��Z���Bye�"�'�|�1�,mW�V��ۡ(/��kl+@y��F�f��+�ύ�|jL>Z�������8I��=��V�=y��㖪��ru���Rؽ��h���(�#�V�/_���r�^�T5�GQ���(�C���4(�4˶b����F�fي,������&9��#9Ɇ�w;�hQ^zy���m�x��Pd�ҡ0�؋bv�n���)��l]i9O����)��Jg�����h��jS��læg6�$m��ms��#�
T��x㨧�4�ZP���pZ�s��|�Ɋ��M��)���i�_��	3�t*��ۯ�.��w��ZS�u�7q��P8]�n���cӪ�	����ȝg�G�H���q2���얭t���|��M������<-���}�`	�cҌ8e�B]7���%p��h�x���0�뜳B���|V��ܱӞ����}���M�-��t���3� �����ڽ�x��2�$�kh�hHǩ��@9�7b��?�p�~/�1_�Ё����'a��}�]�ֺ��c}+�iSf��Όz��v����v�y��1��M\�Z���"Xv��3��>�r�����P��C2pr u�����Z�ߗ��2����ӅD���	J�I�/Ą��2�?A���)�\�9��@|)�F���|X��R��E�
s�<:M���L<�~Ng�]U�/�!T��fg �:�P�&;ڳ�����=�l��N���uon���&U�h�z;������ׇ�"yk�Q�x/aď(<��G��i}#	�+�T��u�w���G{7�lG{7*m�U�h�Z���,+��4xH�w� |P4�Au�q��X�J�=�E���&�/ H�j��ʆ'��!�|�e�p:&�p|L�L�L��9r-c�aE���ēl��@x��|"��uE��aB���Br���N���Q��Ϝ��v�0�L���}��k�;%���c���G�8��saװ#�]�0;�d=�^|@Q ��	�ލ�"�/�K=2�N���(d+`��e�����@����:�2�2.�<ņ�"�نӊOʬ�U��/�$d�44<�h"��R��d��n�]�2e�������*hcmDކ������~��^.C赬Yi�u��i>mڔ	�?�;L~*`\p�&��dA��Z&.�O�ˉ�͐���r[ �d�Ђ%@^?�?lt��kS�k���ؘ|�1��1�Ա>�3��p�<�wD�#����pqM��9*9&�y4�4�����F���|�ʍ����lbH�_t�h�����\���u��A3*ُ�?rq���	4��{�=�#����VbdZ[�����ʈ�1]aP�I��^Ww�X�t4��i�)q���G��k�K�R�� ����:�g� �'�'�)�U9>apd�s�Ѫg�wA{7�iA(�Ґ�PG�M8C�R�s.�R<vYm1�58��_�(�Ȑ(�����ʃ�B ��������K�ڡ���	zc� ^��Dϊ.�Ī+��C��ܫ3����9�~Ww�Q�����bq��s��>^�5�G=�\�Q7;���6R��Z�[w�~<��p\ѷp��j��>���܄:�ߦ����d{fbb����V�i%`,���mů�����
@�p�~�_��{���D�L��=~ٖFT!���a�۷/��_�E��}��v�UW�g��O�|�W��e��~�2 ����)MA>"�t���I�����c{��c���S�q�� ���-B_���tw���>j=�J��O�d�V2�n?M�f� 쑉�'�أz�js�� ��E�8��[�S�5�e�D{e�A�މ���	N.XH�������?}r���"�;���Y4#��y��㔋��u��iZ�p��=��\|�����^��w~XJN��AZ�v��U�X*G�ε,�+X`4��4Ui�����wJ��e���Pbn����ئ�A,"�6���5�S	^Ta�'�:*ζPm����k}u� �� �1n۫@���P;ך|.���y)b�I<�sP���ԩ�ma����� �(j �,o;��ڑ����t�����Wt<����2�T����>��60;��݅����o�� ��@W�^�=��L>��%Q�VR��Y��M�Ϗi��G��${��Hnw>���׎>��F�S����KՏ���C�%�hK�VE�R�!����8����IS���&V~j�'6e�B�� '-�lj��GKV�21I����z����ٺ}�����а�����&�z20����/�3s����M�nR��!��\�r'(l��:����'��ѫh�U��$�'lO'ƽ1�+-~�yL=HQni�#��`Դ�"��u���d�X&o���F;UL@�6P�e����|Z$�(���2�e��X��n3�E��p,'T[�LT|�$J�O�D���f�%_�Jq&M��P�)TD\	��'�W��W�QW�U/o����y���1)2.#��9�Ir"��e���|X!W�P��'7&�r����+1j�6�Ĝ �?�ߢX\c������l{�cQA
=1���Mhk�.�8���>۱c���}��Z��z>�j��x@���ˤ�j�oA�-}<-�9�v0����ٹY�������Ky�C�5�����⡉s�;��۩�U$�PiԳ���7�YG��e� ��m�5��u/$е?�B���R��)�����'ѳ��>�?S�|�5���!s]1�(tu,��i)Ħ"�Օ�V�G���;�t�<�@�����H3p�JL�z\ ɉ���&H9o�J�_>i8�i��FU�� q����[���i�b%�������?��4ߪ{^*�|͢��O��ԎY��&����U�B���N��գ�d��7MS�y}���K��G�1��4�E�Y���%`׍��ZҒ̄�7���j��1��ʴ˿o�c�==��I�R%�L��x��R��W����/�'��g ���?�v�S�Bu�=1��P����ӝ���i����)�Z�T|!��24��<'3�cH|[l,�&A9�A�.[�On�ɟ�[�4"�����Z����	?�R�<�4�TQ5��1� ���yy}E�������$P�f)4V�1Ƚ3	㓏f1B&��M�6(�y��x�d��T
_f��&D���V�o�Q��a	�2��r[�u�u�OI� �]�L���Y�@��O��-c6`���0�j���ޖ���mX��<�3��{&Ս*���}�����$��4q��$�[`��f������Q/:F"��c���.���k=U�Ў`~���A�rF��fp���MA{;����?�Nꝝ�W�U��<�E�ex����ą~��M�ʵ�
�"ŉ�R�	�@���l�e�_<�!�S��pX������.OȒZ�,��¾���\�����N�g<�#:���? ��K9�ޗ��T�oH��C'��@��х0���1`�*OX��!�����&DPb.0ȅJ��
e:�\��2�&�֧t�©��=%�J9RSSlk���@���qo�xN�&$�DEZYG�@VOD��.����?� �Y�����o��%�H���6t@�o
9S$�+��Kh�ď�cA�k�W�oې�r禐��		�A��U��t�w���颮�d�Uh�Ǘ ���	���Zv=|I�	�3�q􋐰A�D?��~�����+����F�v�_#Be�"^�RRf�q�Y��h� Aɇ��
��v\
��ʽ4�M�	 eSl���IF���8x�M��k���X�{P9R�f�LP���g��8du�Ը�E�l��G�J���ŷhBw ΐ�@�Ur��dk��\'bP&��:ʕ�!3� ������=��@	vf�\pe<p���F��R��NFzYg��W��9E;@���#��r�~⦲z%-'3؃ f��ݰ���Zu��a�s��^7�8�g����>X�&�$��,�Ov�v�]�Y�����I�w�֮_c���;��>e2����U=�Y�5�Z+�.���'��xf�ܹ�I�m���W���1�`��e�24��|�=��>�xx�o���������(m��Q:6B��ز��G6��s}6�3��tA
-d�?$���f?GE�����Sr��<��	~%B�7@D
��<24eY��r��]Dz��/�˷B�?�Y�3�s�5>��FN	x�����A��B!N�;B�`U���;Uă�d�;;a(�i�t?G^�v1削c5:�k���xHsP:]�aND_3����M�K8�A��U�:�qSTg���~ޖ��'d��u��TAY�ML�mЩ�S)�	zS��M�˵���*��A)log�U@�B�3۬ϊa{n�	�3�Mbߢ�	�lMN)zD�ܯ������3��S�i��flnv�-�	fzf\46��kjb�jZ��U{l����ҡQ�ȝ�����FcF�,�9�x�t׽���v<.����kGlhh�} i��g�lnF}13���O���?�>����y!�<�����x�B�rY���W���څ$ה#?�ϥ�ϼ�[�Qԏ,�(���/v�`Q'OS�N@��/���m��Wȣ��`��3ǸM�l��Li¥LAf�����3dAT��"P���'E��
R�Q2�SAv�:@�8V��ܕ)�dp]�xW������5�l��2��r�	)�X��38-V{mq`�u��Jߐ�L�ybaZzj)�ML!��v�Z;x��xw��� bĵ�nY/��s�@Y~�rD�� O�Ej�EB�t��'%z9r��8T%Gn6��!��B��
��8ϖ*2d^y��&xF���T(�O����B��;T�4�|��Q�%k�&�E�����gm�+��y�S�k[!�P��A���z�$_�����B(yz����r�m,�+�'L�Y �&��n�`�A;���Zֳd}�=V��F��x��ܕ?X�X�I���O������ŁH�a5J�=��|ʜ���ܩ����.oc=�>���G��m�沤�6��o"}�t�]ݱ��{9?����kN�C���Ǚ��x�NP�E���ݕ�u�Zpߗ��9�6�(<O>�蕐A��D��:��*����t`��>o!�%ŏ��αE0���� ����Q��Ӧ׏X�S�'�H%��	.����)��7c!��j��[��W	FoH'+�m��/��ϑ'g���_	�����������D���k�x6Ņ|�mA;���[���e�ߗkڤ�t0�h/O(5��8P~���4�:�
���k3PW�^��"ߗ*��p2�r?�h=؄����A����1�\O���w{��2��l�~�~����v��[�~�~'�?>@D�ȦS;r}d��U��IL�v����b��_�sD�֕��P�O��#��T�y�G�/�J��K��	�t�'"E1X��ea0+���T�R{�,�.: % ���hcgc�����%r�><]��e�M�̋$1c+�^I�eu�#����>��x��͉4M��$�>(r~v8K�q�	x�/ e�S��Τ�R���)a%p�$�"��U�;|}FGG}�'�q����D �(��Om�ޑh�W.5�� I�'��"�H[5�}Z&�v��tΧ�յ.��B<ѥFC�P��:��J^�<8���\��\0��9W6u��2x�2���l�'/�)�0T2���� f8a�?������Z���M>�
<!ES�4��)�"nO�"{�9���KD\Վ�;6���xH|�ްaC�@;�i�@Z��[�e�|�A��s"@o�p o���D�d[ڱ<4h�e9�H�6GS�f����)L/}���%l�ԃי�#�~����>�8�����v�Qr��=m\�Ԑ��Òp��f�P�<R�/�2-��8[w_�ELGz΂kVe"�$4����@N���9�����[�v��+ms��]f�=lO����,�7RS��ۚ��$����ԇ$d��Bg]�ӛ�2���Vc��(����=�5B� �
�k㋄<~�/��L���rˑ/%uOe:� �G+���������i��xz��D��-��-���;Y� ���\�r{N�m����Çm箝�f�F���p��}�f|�ߺ� >ȏ_ʃ9��I���#�8�v�6ƛ/R����� ����_��[J#OQ�qv2�\�.(���(�N�-!w�7FeV_�(U[v���X�)�!�P*I9�?�HQ���KZ�����(�Z�B��d ����<�J�R,�	���*P�LtE�gQN��
HB���T4:խJ�^SR+�����ۡC��o����?�K�z��)�������M)5�v�P��5�ɒO��e�@�r���vB�mLҀ���r�JƔ�9�8���q����t��i%nQU�jR'ՉC|
@-%@v�HY�:3.��
�0KՖ!f�V��r�W^��5�Ϡ��
йapAǴY�!D�C'>'K[�@���j�uzc;=
�A���C�~؆bɮ�Z=��$/�k�'����͂.c��6'&1"q]�*����	h%=�GCҾD�O�>��wU�Ə������O��!��ʜMȟY,ے��'T}�?�C�*5��z��8ωW��.=O��V�W�b�R�&K��'P�a�x�"�f��i�pԜ���.J(�_B {D�➦��W�c�!:�v����/��
��+θ<����{���ְ���.60��HZt@>����y`�+����@�O:��rJ����N(�;t��T�ˈCI�I��$@��0�1K�{j2�J����4`' �9�E� �J¾���d�.��1�[~���"�X��vt�󶄝�H����-W��]�3󽟣�G�Q�/e������&'&�鶭[����P聾�E�C�U��}N8�y�d ���r�w�EQ�b�6 �L���.������_$��)�.�pL$�A�$t[vUDz���NhKC���[��Y�����4Wm؜���Q^u*�7v.,���>��7������,�@c�I��$(�zHb-)��Y��,Mu	���(Ol��tV�C���%�[	���;��t�L��p|���~P�-x*�M�]�P�OL���+�6T��J;*�Y(�(�w;d�NC.R�K_B��z[@Y����e� �{@��W����u�H��k2N�_������ƍm�;+t|����Uʿ�_���i�o	��K�a#��RS}n&^~<���V�И���1��Z���7mSV�ׄ�`kf���X5ĩn��Q��^�Pz)Q����yUȂ>d�?{զ�Z�dKk�6ԘR�Y����Ŏ��K�vO���)�W`��fM��1��ފd�S3ƭ�RS�'�,t�m���/�?�&Z�ס���X51���j)�V�AW$
�_�_3f�$'@��5�����%V��̮#$a ���)�${E�osH*j�A��W��/�� rU�id��繭�E�=�ek�HЌ��EiE�2_,d�#,[�:����6�k|��O_9�Ϸ4�j�O�s������>���4`K��>'!S�I@9�³�*_4����:ڵ�rrQ���w����}��y���~��ϳ�#��v�_k?�����8ۡv��+�o�}�r䚈����x����4M�ZmB^��g۫������+ֱ�a^��]������˞ko������W�#6���?�`�"���?��ꍯ��}�3l�l�Ff��ig�f��ϱ�{�3�w_r����smm��.��/��zP���)]�4�AOFc�eܩ�`�����> ^��"�L�<��2��Z��߷�ZxYG�u��&���u*��z�*�Kdk���.�D�˴�%�ɳ@	��D~��Ҷ���)���YS��6�r���)�T��p���|�	:�d��� \a��;�����H��n��f�����(����[��'~P)���U�&�_��rO����L�؁�ǐ�۫�П, 2r_�A�����<��=I²?��h_Y��J��
b׮]�=����G�i���]����]}����[�qV���Y�c��tf���]~�����gq¶i�z��;��[��N��u�J��f�ɳ�E�:���ٵ�~�O���M��*ꚶ��2;k`�F���[c�����N���þ��=���δG�}�&��պz����!|�C�/}\���Z��� ����8`k'g>%𞢃�yI>qi�����	�p��J��Zl|�*�w���j FS�7	������������>-�y=�(v�A��xh]\@�'�@�x�;'Ͷ���c ���E��due�������:����aG|�g���6('�m�6� �>�'� ��>$E\>I���]�]nc�/�Kñ`���H��#?���7�Ŀ���@��ɞ�|�vD��������i�����FlK�]v���^��Flú-�%��5=��w�-p�=�.;{�z{�������g��_���k�ڱI��$S�&�9���e�m�l]���{���5��u����S����n{��>dz�m�w�f{jֈg
�ϖ.�C�PnP�j��elE���983��,3/іg��97��N:Q(ʗ�d���_��?�N�kWj�;��c->�m�9�q��Ԅ�y���a��O`��0�p;f�P�er@��Aت;L}�$��"�h�Co��e��и=rԿ�w���hڸo�>Ѥ�ys,f�̓�'���u�^�t�0�,r�>�|�	[����M�Ia�գ��J���i���ɨnC���X�R���E����cV��:M@瞿GܺmHx��3m����Du��Us��=#��:s�:[g���w�o_:ذ����[ߺ��ݾ֦�ݶ{]���㯲��ñ�u�K�����9;7��#vױ)���I��ȼU$x�d
���"��vS��ep�b
�����6:�FV +;5J�/��R�e���w,W
�gl��Q�#�TƓJƊG�<��ZijuY�ז�KD�V8�$�qA�V��&��UgZ���|w��@�����:���L�	���<�Kz<}�������n�j����= ^��dQ�͠iC�ɻ;��@�{w���:��������y��F<��(vCMQ.�v�b(Nf���<k�Ex�c/��>���+ϱ����v�ju��<hC���{�]p�.���-j{r��ݶU�GO_����^q�I����a##U�T���5�C:xdƦj۸f�K��^q����M���)M.��*9���֍�kG�����/��|��H��Ơ�SҮ��Wz�������YI��+��#|R��(�:�0D���p,>t�:�����a�@�:@��y%k+�����2��X����J(ڱ
<q�R�2�C~����S�O�^�Nr�Pv@��c7�r͛/���>A��L�d}�c;@�:f�
�z(S6�NN�>������=�ۻw����"~{A��V�������}���ѣ���g&���N�p Z��_c��b�I��M��:�a^���ID���?jq$^��=���]i�������X[��g}ܾ��u0��%;�������;z�=��uv����[���[����h���وv=���h���M̛�,V�6c�1��3���m�Z������XCc��k}�~�ܾ�z5�m��˷m��y���[�}rX����c�J�I��wxJ@�����v��B�L#:�dr������n�Dټ�,��&}�3���ݑ�(���K��8M�� �z5B�&�x���V��\������a��8��沀�2���V��C|W��5��@m���I��֎��,Gb�6�R��@uj@Po�<��DD̏V#-�H�K���i��9Ȓ�c�H���.��ݕn[�a�?z<1>aG��.4���V�Ԧ���;<�k׮]~�x{��4=!����=�?�@J������6C���v:��sI����>�I)<)���cfՇ���v��n���p���7��ɧ����c��sN�M��v�}�aM>;6��swn���X��]I�^|�n{�s.�����]ۭ���Ԓ�Z���^�|���-���\��v��d�ߵ_���XUuUD��D�X�O߾���ػ>�yMj���G^�u����vG�ڀ�������A�-)\;cE4���g��ƈs:�m��ssn ���t�hU_э�n�ɤ#8}B�(�����!9�6h/�<d�iY>�eڇіV��@��T���0� @����b�2���V\�}�%��SE�@�ގ'
^�$Ka�E�)�?��4�$��ݑV���c�4�0��Y�	J���������ět�:�(Y^��X���g��'B�'�-m����[�y��ɓǨ9fc�����.�L�|]`'(�SO;������.�Z��l�� ��١��\�B����nt�ڽO˧&�@� � �=9_����{�������ݎ��ZC;\�Tm��c65>g{v��y�၃v�q����ܰY��a�NMeў{����'^`�鉏�Ӵ@���W{�l�v@L��6������p��y0�L�ͻw{9�pȑ A $@b�EJ��l��m�EY�2?I�,YV�eˢD��$%�@��D��pw���6O��?OU�;������dv�Լ��������4�-��^��,w���'��Z����]q�%�p�у��?�[���į�y?��?�=�7�\��T{�{���c���WBD3fAN#Њ���\`e��W<��5q����`�2��\���<;���K���F�x3�d�L|�SC�3�Ep	�&������Na+�i��u��	�Ac������j\B۬���%��Mv��׸!�pD�#N�Si	*��|!��T���׹��Š�<W~F'�՞�k#�_���j����9���������5����y�v�ja~��}����<�B��H�vgWԫ�Cy�w?*�gwt]GS}�c�{�Ge���"4�D���{����r��*���Hq�6<_��I����V��-��N7�GRRVii���T��&rZ���)d�h�86u
��
:�G��ɩyhɧ'{�{��T8�2��{��}�^��_߃G�Ǒ�
N���B1[ǖ]�/�@�V��0��m�y[�����p�𢍓8��W��@.x�m���}ܿ@0P;�G�T���s��C{G�hx:U��+����ہR�8{�^]�6�ӛ�Q�)����f Aɧd�J.�Z�� V�:h����9RF��`Pvy�U*A�"�?e�a-��������p�x,o<��'Va�/F�A�]H�6�-��	�L~�\u��٩>Y�i��=QN���Il�r����	l��+��r�`@�d��#�]m�(*��S��H����D�^��с���=��`|�b�8��t��o���nI��A�$'�;�t������ ��:����ި�낦NNa��b�%��_i֋��=/PQ�x�mK�[!����P?�?���PF�X���)^ ��ӁD�ܺ��V+�c�0����F%+ь)� �[���v��G��G*�8�,ٵ1�����x��QX�ʝ�3�Np7\D=;��>�(~����>�8^��S˨W[xݥ�Gn�?|�M�Y���9�g���g�i���(~�S_��b���Ǐ�G^�Z��7ގ��-����:lg=��	��jl���/����~ә�bl�u�uT�C��JA��*��C5��O]��;]�/�-#�c���C��\�-��P��`JT��G �"*Oz�c/D�aA�)9z��#A�`�t1,�o��4�h�w0��P�n(Dk��z�-��#�j��y4�I�b��T9,�)�4�)OC2I�[��`M`}f�Ԧ4F9 �.�jkgO��w^2]�̡xh=1�P��B�������
��t�FFF̠KE�xr�]j6����i^|D������-?��:�n&Щ�cG�����Ilۺ�v;�_�������೓Л�&�R(+�������n�Ɓ��3vU�gH�Z�h���Dux=iP�?��F�N��Ȣ��s~�_�׳E{;�^���4P��`fQa?>y|ӕ�y�(N��8�<�c'g���Q�w��|�s]O�d
�=;�m�#��oy	.�܈'O��S+��ᓸ��%|~�wO�Xi`ax�p�~�	m(�=�]���xf�j��G�χ��-P#�ܮ�l�0mT�����<qbu�S���0�;��
��a�t%)�hr@*���3��๊�tOQ���p�({�[7/�7�2
��c��-�����l	����u�fbr7*�!]���=���@/��P��t�R�JӃez[��f�v\󔙼TD�G����\9�kq��� �ce�N�����&ob^��9�W��TGs@��{ې����W���2�w�H6##Q�-�>v;�Jj���D�㌨}^<��#����AT	�W��e�Z�x�!�[����h���hrxy��&����4��ǴR�aǊ�>�'Z��.�:M{o�9-��nH��%���i-][�.HG�����M�g���术z�.��n�+t��W��7�L~�|�'ʤ�!��$=��4��O8h��U_ȭ��<���m���|J�Q���xNU/��v:cϏu&��ȣ�h�cO��<r-� <;s
�>�Zc��qtjx���?�D*�j�k�kvp�#p����m��cx�ٓ�o�Pj�k^�L�vQ�L_{�.ۘ[�s5��v�ph��>+p�����vtZ����G�����>���E��<�����;���O�b�6Gs9�����Hmj�ά���=�t�82�V���>�����skY� ��p�:h:���EÄX?i�zT`�ޜ��59�'qR�	,ϧ�Ejw����5z�����c�� X�@:�6|�wW��NRe�b?ƿ������@ �;y\p�͘)oB��nљ����	1����A+���;��A��
P���6;����9rZ��P���r*����z�J��D��B��"�jP�XnT�ד��up@��8�mcW�Cz��Xj4q�Fg��Q��]h�X�<z].A��q�W.����w/�&
)��8TB�0�J�I��}�L2D	��T��J��ejR����J�#�O��h.�P�|�r�C}tؔ��J�Xb�Y����Bۅ���p^��8n�7`;h؊�i<��?���i��]Ǌ�*e��Ġ?%��(��ڈ�)�г��ϯd�2��l�w�{0�5s��L��*V�uh0>k@Bs�FH�;[P�u7\��@�Z������c�sA�<Sc��'Dâ�D�JnrE��98{ 1��l�<`Q�{;��s�X��$O"[�7��#�o��7���`��Q��Y��I�CCiԅ��A��6`�n���Q�,�7t.-H�4�y@r����=�p�T͈4��,r�V���,�����B+�1ƱJ��ϔ̞�*U,)��E�eKt6r&;���s�wB-�
M���V��e���,9�|�T�u�#5�
�m��KvVzFe�읞BR��zSC�S���������C�?ۻ����<��b=����@,?�T�#><b����(�L�)�X��[�E=�L�%X4=(tԊ]-��@(nr��R6l�ͭ.��#��'m0	��M�u[���w]�W^6��K9<7=���?��r���-�V.�q��l��{���rn�hW��6��?}�>���.���,s�ȫ.���lvNdq��sՒ�`�`��w]�?�-��W��[o݉w^�[F�RZh�	�����I��/�)f��k7�'^��]8��SM<�2�B~���㽷\�͛�x��u\�-�W��o~赛�֗��%�F07;��e�4�.o�t �����^�ox�n�ےŉ�
fVt{f�|c(���z1�y�N�,Wq��D�K�GJV���5����m���i,c��#��a��I`�I��Mx�-A�Iԉ�8�(1�v���
��b@tz��v>���2TV���k`Һp8��;K0�e��z9���s
�)�C.��rP�z�+�9,��嬚\�4�`���Mz������-�[k�Ho'B�H�9����7i}D��|�oS{U�S����ꃓh�mC�<l,_~�ò��	��>U�Q�zu�������2\.��I��ѵ&ngۅ�;��1F�աh��]�cZ�qy����=��2�U�j�^��EG[��irq�[����P}���'h}�d=:�.�՘悊K^,�?���/�,�J��=�y���[x����|�$%Y�AQ����&<[Єe�4i����Z �Ld���c���bj���N��3�NOMiY�ѨY}MKG�8��	�e�=y��|`�8;�F�
�ߕ��;p��Qt����6�Zx��2^��@�QƖ�^z^7���qM��l����]\�q �l���g��o����=�nG:+�a�5���d~�W�[��0�f�+�Dp�ة/�����Y��Q������@߆��o��t�<r(Ӡ\�m��;^��vsGG6Ti���G���t1n�>�a,��6��p5�ؔ�@��	N���ۈ�|���3�y������]øuwW�oFI��R0�la\T���a�4���Yk�guR+@6FG]�����ʑ��;��'��q�	���씤�-�!��n�a�&�<圪4�xu��L9�8Nut����ֵ��9�Ӏ�.��%s7l�;�t�E�Cu�NNF�P��촙9���8�Y�lʥ2F�k�8����Mm�S~��5�SS����F��]&�~�9���=X*N����n�o�nb�\A
��Yt)���]�):t�t*Ef49��
�����N{��P6�څZظr�
��9���vYt(-��r�b��ǢݑHR�#_?r�i�t��AC
d�=?r�kiJ�������$�(����
G�{A���f��ZEhI~!�s5�#1���2�Y��P����<.�
��9	��*ǯ�&W���zŸn~P�K-��9j��:�*��`-��~��z�+:V�k����^�A���DU���ڮvP�Ž~�N��=xd�l3�m�
��"Vt6�y�����/�u�`�����A|�?�w����O��ؿ0�k7v���؎���+1(R�+Q�*�i��A}�>�_��'�7����u������[�Q�L:�7�z�|��d��qx�������8>��K'�xÍ�}����\0�?Q����g�+��oP�,㪭C���q��:�]��{��\AQ�Y���p�K!']�)���t��n��cG�1��0�*�w��?��	2�-'�Q5�CY;��2����|�M�B�+C]��,�d�&�ـ�e~��ߙ�yz��$6�©1999!��������Y"�b,>6n811a���o]W�v�I���h	� ���6�e_8H�\6G6��a7��ch���d�bT@�X�gсD4{p����hU,�Aj!�6m=w$�$ك8F�߀���I���ik_g}�4��D0.�C��qH�y��"2���y��?F�	d��[����wo}kUaB�ֵȣ��)!(� �$���N(��CT�r�ڮ�@X�&t�Rg��b��dWrRR�t/a�|EH�+Cb�cM2~����LW�he�rt4��3;I�b���/ފΟ�A�;�z�z�Q|��4��/6�ÿ� �9����Q��cDF�`�)j�2V2���O>���`��{�e���W����&�n�z��ǎ/�3e�5���w?e���][�?�����?�~bw5��OUq��%���k�c،����2��SrJ�!��$	�.A�T�Ky��q�R3N麖A'#Y5�̙0ͯC�O��,��U�&_@��<�2~D=��Q����fT��kg�O��:�%�XU?+i���Oիx�љ��1�xL0���<���P����S,�\Pن�ƽX,Mr��9}�K��.Q,��3����k���q�~R52('�y�0_��C$�ȟ��5ʹ9;����h�`GP�-�BR���e<t��**�xx;9�Oˏ"��6`R�V�>��
z���-�L\Y���ߴ#�P����S|�Nd9�⺼.��]y;�K�A֯��d7�(��j�.�Kf��*��!���/���D�<�/=�w?Z�61�]���O���_~��tp��A�?�U�_gf��"9a�.e����*n���f���g���M����*Mby��s�6V.`�hN���r��cKԸb���c96u�@���6E���mU�ճ�-�i�P׃h�h��:W-'�����=7�r�f(c�a�d��)	��1��|�i�+x���R�'k���`�Y�;\[h�\R��g�����`��N���(�Bi�>�SN�����1l���*`��'�����}�s�����:����G;���֔֞�g����te�s���4�ز�����smS�#,ܽ�5�{Au$����6!PF���D�ƀGu�MUH��z��c���XW�����΃掖Sw<	TO�;(B&E��M"O@�ʒ���Z�Hc�mYe0�O��+���S+�r�t��gY�3V= �=H]荷�ZZ����B����r��^���D��R�K\�w���z)+*r5��6i��H���{�@c�C����Jظ��7x�x�j;�R���c�.���Kt*�_ѭ�� ������S7�e�Ch����;�nyمt$y��<�?w��(�kgF��Hsv{f�u� �F�LJK(�Xa��y����Ҟi��+�ư]���z�Zm�y�*P���`!w�XR�4�~z��mc�ǫ]����c7����Hk9|9 :�<LFwY]o���Q5[�T����&w��;;8�3v�W�M�.�$'!���s�f�F�N�+~s�
�#D{�t��Gi:C��P��j拨O�1���0�F�yU�P��.??5ϲ,��qQ&���s��f��괫�"k��q>�M�[��FtI-��r�� {�������zQ�ȋ}Hy���(��a�.���}?�%�[m	�u04�YR��K� ){�(�B�R��<M��6�> ����X[O�kʰh r"X}��z�B6Q�]��L����2+t$܉ܾso�d�}�&lҫ3
ؾ��w��ۯ߆�\D�8`�tvz�fi�M�V�=�x���}7o��u��mN�]������T��JP礪c����[�4�&��hkstJ{6�R��r��-7o�w^��z��oƣ���B�.���d#G]�Q�jE���k'��?�&���x�L�A�9�Z4���*̉��b�Ӷ ��*/ԇ�4F���&��}|���T�b�IGa�آÑC�4]��SѮGƆi���\�PD��՝E���բ�m�r'9So�8�P�}ܢ��輥Q��G3֒2ն֎5>gϗ�e`��x�;�Q�J����	�lޅ���C�~����Ϲj,m��֮�S�sϋ�C��΁�i��O"ԙyGZZ	4�1��J��2�� 6�_�Z����XZ�j�׍OBbd�6�q=�FΌ��eP���C_?��˯�/}������Gc���]����_���f6ۊ�u�ص�M<:��/�G����d��޴��v���m�vK�SGO٭��o߄ђv]EԸ3�g�t�\�g�p��	���Hg�ffPj��j��v;R���W��޸��?��,���t���专1�C��N'�M���p7TF��Jg2����h����
��&FF��i���Uq�ďƛ�9-��An�M' �K͆6�B8`��/��dyB�
9� Z]���
�D�h�1���8D�|�?���F(���t2:�&�c��Z9ҋ�;Z{Kp�r�k�tr%:�Np�p�;�F��; ���G��]J[�Xe|�^4l>��Ҟ�a��� j��P��EؠY@?�Mn����ΐl�l/(��I�@i��g��]�P���?{8�>�k�7���T��f2
������3+D[�Ӂ8�-�<ƁmN2U��bс��[E��vI͈�m��|[ˍ��T��r��P(���~��i<|����4>t��x��ݏ�����<����=z�����g����)�Ȭ`�5�_��g��_;�Gf��?����#���#t*4�zF!��<r�4rWm�K/+a�TG�]�R4��l��J�<��{�����\	�]l�D���رe��pO������s�X���,��mkhD+-�X�q�6��#:���Z�h[�l��p�7תa�vx������f\��8>OV夗����CY�Jt��ө/u���Nr]�>�a���m����ˮ%�3	G��_3M�#�vj���^��]cF��3]͵1��l,::%:�l�@���'O_S��b�rt8J�����Y��f�tBu�W��^���C�����@l�?4�Y��ߨ��L=�D�uչ��nGs�B�~&)Ǘ��S`�2��
3���1T��_�� 9�Z��q�v�	Wdh�A��\���K2j w�~c��6?bM������C��-6l�G�<����N�����m�u�2���F����r�=D�Z���#M���O7�M�0X��R��ȇC��cb�.���Y����XcRTr4�e|������#����_�'��3���#���N����|�#���GplX)�P�q�#'�:�?���9��mW�������e̜���ce��4��v�brZY���2n�t~�%�p��2��Y��g�'9��no���<w4_}`?���Y|��
��ʙ
�p�&�,�:��}���vg�0w;�+U���M7��d)����§�{
�v����%���|l7_8��^9��v���y�shV7��ae񮛶`�����J���(���	�S���G\�a"�r0
���UkUp��3,]�Br *&��(�v��DG�zs]���V���G���~>�c��u�NN�4L�m�v�5�y�m�8oL
$`R�>?O�3Ȗwf/8H�\����M{�/���l3��/u���⬏mEu|���\������e>
<#����	��3&�Jwë��L����Hz��I�%W�sz@<B����t���M[�K'���pL1�l��H�u*��W_�'<d Mg�]��K��~��#z\<4�L��1C���'�L|�� z�t�̡��<�u���R��k���W���x<1V�V�0NZ$#�^�M%l�� ��eiNp�s-5N��L	G�y��h��M��n�Xa�� '���Z�|}K�a�;�(5�Po�������~�c�p������m���w~�W�_�~��;��N��ß�]O,�ٮ�\Ǻ(�B�z2�+�!�fG�Z�� ��%W�ҪvH�"���gqba{�s��7���y�y�`"�#K�������	�F�;���{��G_{6p�������8j���)_�:U�q�����/�9�vk��c���z��G�99�p�Mh��)b���	w6��OtJN��|���?���P;�������h((?�kC��b��_�p'�S����{��) �U�Q�9C�����؅4����&=���.����b���f�C}H��s�X��{���p���ۀ��f:!��g�cm�h�*e�k=�S�� �#��->R�3'}HﺜoX]$�ٍ�яN��P]��r��#D���,D9-�~�����'���<�IT0�&��Z�U�]T�´��,?�<�f��,˘�؍��.b��*�@�e�47'ʱ�	�+�S(_��&)y*Ut�Mda�S�c\Ƞ����i����r+��]`�&6�D����,[�*a�^�'�@9ҟ��VB��Wɻ�<�ӄ!��5KG��if�4� 2.iu��`~�^<��#<~b	_��V�����]��Qk�}��je	'���ǧ�+{�}v-?{���~�C~��dt#st:����*^�ow&Y<q��{�\ı��~�&Ɗ�`;VjY<�\��7�G0�	���z��"iFi���������y�:Q�r^�*��u��1�T�ɹ<��>��gq�E�O9�l��!�@wrK��ZЌ�:W�G��MU��N�UNGmTi�)l��y�>$�5S�~�@�#[�<�^��wN挴PQ�a������ޓ�ϊ^׊��W>�T�|�2���Q.EM��&=c���G��T��+�C;|�ߥ����.��T�)������-�i�#�
me��/:�N?*�O<2�4
���e��ܰ�P�2�.�_��-����n����7T��I��gY�ƣ�)��1#B�Z�Me�5?��t#֬�t"�����x�0�YV�hOc���z,]���¢�"���>��6��R�ƅ��f �#A�wI+[,���p���8>tT���̓��f�ʳ#��1��|2�v�^,�}��q��e;oY��Q�zB[�Qqۥ�V6�H ��P�B4L�>��J#zq����Qĵ۝cîW����jI��R_Ԥ�2[�U����n���8Ȱ�tu���A4m:�����6��J\��3DHp^����N_U��z��g WÞ����5�28������$\�-�Ml)b+W�9:�:��J����/� [$
T�z�i�w�����<Jm�V+`$_�b5�Ë�Xb���^�b� �Ε0S�i;��U��:�Җ:l,ccp�����t#���*�Fj��*��ҡ�<n˅Q̷����;5ʦI� 3E����S�ǐm�£_�4
�Y����R���1aE�
|�(?B�§�"�՘�I@ibQe[�Yc�q�J5��1^�0�ы�u�zwL�4ؘ$��'�kLX�o�$
ё�Q8�[�r�y�HK�յta�&���2B�y$o3tV��{y�ٟ.e�����N�4 �����eD:U9�����T���#Z\$���Ł��z�ڝ�G��.W��B�$�K=h�:��8%�R�9�Ӎ����ό�΍�H�2���c1�[�/�Fe-`�X��Q��c���b�>K� K:Y`�0��|V�/�;�0|���Ţ���~:�fp>�H��K�"�ש�$��H �
����"�c�X�Q�9�.�34l<�N� 8�]�'C3?���8��o��xD9�@���$'�UA3��ˊ����M�z��M�-m���:�!��q)� =�I���s�U�P���h`��V�|_��{+|�qV'M�!˕��ހmʍ
u*����8 s9�Na 5�9�^a��P�
_
'�:-��l�n���f����K������O��������L�+B��&�K�\bzc�^�Y��Կ%�ukv���4I����SA�g��qd�x�k�Bs��;c�[�Ѩ{�XY�3�[�*우߮�����M�=�ae<n���������`�D�ޙ'ARi�.�Ԅ1�Z=h�4�Ҹ��t��.���t��t[y�cm
1��W8-?�������e)	w .�؄r�l�2��۩躍wv�T���_;�h˹�B��Y$�P����Ȃ�ah�"��Nsl��(I")d2n:Gj��� Y&Eg���*�X����ú������u+r]���g��{�[���Q(����w��܍%�6>��	0����U��,�n㜕������y��}ΧQ*���]njp�/*ʳ	k�MZ~%���%[	�W��g�S	��9Ҫ��&M`⯴�4S}pfNGGd�n�Dhe)��'q�`=��|a��e�R��i�?�>�ߜ��8U��@�]_��B�;�i��k�в�R���kF�@��Qj�3A
뙰4Nz��!������ajR $�.�J����.�S�:'�v42:E�
���K#�R�Q�9�j�t�y�Ӕч�>�YF�tZ��-��p���lu-��'���Y���0)^��KwMN �O�1k�酌ZPi��BF�i�o(.Y��W�Kh�E�0=���h��U��"�B����w��ON繼��9
�">�H������ꫜ�FKs���>�gsP���d�u8'0�#�n���Z�h��ksr
avBs�<�c�j��B�X�ʄL�	�H��,�YȰ�A"����2�C��f�nK�/��l59**�y���|��YҹXݴ�,�n�_�N�2{[��N���'�ȍa?E2��N�f!���U�3�|��
o�lO�������K�P��ܪٟa58Y�F�Zu�b�̠%��;�����0�OBX�wH����R�:�1�M+���I9������$�ă��9�*;P����-�Mz�Q�nL��ЫN�곮O��&�o�·5%=��
�!k��C�������������2يKze��[�z�v��v8�VH���{'�Rt�J�Go}�h�"�>){��^���Vr��`d�N�J��"r230���j!�ڱٟX�F�Pu���q`�X�A���NE�8�����G���Ƚ��R�O�e�s�&�|�M�K���XY�(]�De�Del�2&�ͣ>6����Wj�>-�$�<Vn}�p�����7
���F�@zJ�D
�c�>�W��V^d�+=��/ȫ.�ǽ�b�e���4�LFR
�ݎhrDtga�\e��ǓUB�Y���R��ıj�/By98��
��dU�O�����'}�/t�(7�8&W�,�x�x�\�;�6x���tfٲ}<j�n�`<K��߬iI��R�(���� �V���nq.�P�3U�1.�˜kM�ڻ_�o�l7�Ap>�K��6Tp��q�Vhp�45���`a���Α���A>'���yo��Q��4O�Alw��i��T�
�:k|B�T���O̘�* E4���|s��ʏ�NE�|֮n���j�Џ��-a���'M����׿q��hƉ`�P�Q�R4��zH2h9Q�lv^H�G�5��ge���T}*h=D�AzFu�@�)-�Q�0C�u�"�M�j串JW~���eM.����]L�j
��M^���8����W�t�Ѱ�)ָ��3�|�0��v��SM5j��h*��>�
����C�#1L3�:��O"5C�\u����ʉF;R���2�'�g<�
������˅j\7�L
��B8��
�4�Y��3O����a��b	cD���TX�2�2����+k����X���I�D:��c���(�AǖfyV��5��[�Q��3Zk��)�bX�F+٬��ii��X��6.���)��8@��!���<8JF9g�"�
���iq��S�}�(p����n[0�zMN}D�v�vXĲW��YI�ˎ�lF3W�Ja�w�Ti�m~���u�b���,Z��5-+l�
C�L�V�3 tm�{�^Z�(
��K���ӕ��[˔�0:�+H�?c�h2u�"]8�X�m�u$�U���}�w��!�)G@�qROڇ��,)�969HyT9��.�ܮڪS>�/6�JiɀG����$C�e�*��Q�W�Q�C]ah�A��O�/6 )��d����SR�Z�k�����o`�m���t/F0���6�F��S|Ic��ds��A��X�����>e@�s���6��j7>�u��y�DO�)?
����N����z��-�~c<���~4��.��� �c���j��)G�����:T֏��:/�[��1�[]�e���♠��b/�P��Ѯ��S��ی�-%���*yY8	{��k�N��u�/�a���m�q�㚙�f���<ǭ���G=�k�"��\��4ԫc2���q���ҿ�}
�������8۫VG;��v�z�N
ma��L��~����בȣ��N�2�\Oy�[�E��ۘ�����&D�2�X�n2��5�v���c�Ł���f�V�f������(�ltDѵ�n�i��C�h��Q��}��Z�r=Ly[j��y*ӑ���M� ���
*6��Ay1� �U��<��(/�M �dk��:��FL*�.�!���ـ ����k�F�ق��=B� ���Z#
��t[!�B�/z�ׇ��IH��4dܧ�����t�����C�{3f!5)g�4t�-��>ZX��ө���[=�L��SO�t$�.��Z,�䧌l#�9!���r�aW=���)ϛ����0Z�D��Fɰ:�y��,r������&�]��;�@�\Ĳ��;��2����G�OΆ��h�ZL�i]��θ�'�2�S�Q��������J�@Ǯ3b܋��ư@rj����ƹ�� %��� �6&��Oi)�3ʪW�j�\�^��!��!���g���@�M�y���X_k̇t��������V	��4���nL�3���.�G�#���`DF�w�j��Yk 1�ʻ�2�Ҕ銋aa�j���ئ�AK=xv&��<N8���.ҽG�PO�Gg7�h4N2�~�����m}.�F&wW׽(#�;��ɧٕ��-é<�N�)��� �n��/��f�^�����8i=�1Ș��Lo�;�.��D�?�#M:ϋ<�-����M���9���Y&G��v�%�!O��g��*h�/V��#�p��GŻ�F0|�>ޟ��`c@	��d���U9� "�̸`��Ɩ���i��Q���VA���bb��Q�r�<0�F<3�s�X��y<�����r8�ܟMz��.HA+�f"(n#�b��Nk I�Ç}�:�q/x;\�P��=+K�,!Em��T����q���S�ΗJ��Ӂթ�B�VmR7�L��_9!�i�x����'(h=�D�i�2㝕�oES��Ń�[�ȭ�xJ-Ic8���5Je�wn�uʈF5W`�v�iU�q�t+G�U�3zoCO�����qs���ݙ���`�U>UWҎ�4(��*��xJ�0��.+#�����=�O���v�r2r69�y4'Ű�P�4� �]G�ۇU�P?&�䔤y�$=o��gT�(�H�Aź)6��r]H��<�K���t��N��1���	:i�h����L������*�?��xn��XZ�<U�Aפ���rcw��+p�p�
����&P]R����8x��􍂝F�:C9��2KQ�Hl�%�u��F`�� ��T�g��?*�ސ��b�"����3@f�d4u����-Yb�câ��n��DC�I<҈���}���`|e��C�N@��dTe��l��=�ix��t�i�yT=�zU���q�e����_�3?��a��C�ѹ�~ڍ�`}�?��$�O�y]�1���[��ؐe^�[��az"�����)<{��d��ǾF��|���5�x��N#�0Q;g�@_�� �͓���j�>NNl��,=�{a�u`=޽,֮����p5Ous0�qH0�&a3�ݰ���!��L�~�.��d�..]�V�0�qX���������8�B���{Sp�䫀���w��Ia|-��lpZ�����>M���o2H�~<-�]�M�Nq�
�_��2�Ҝz&71G=���Z�N�׿��ߌ�B�i
N �hLL�#�?n�ϣ�LN};�턭���NȰ�G��w(0qRF��&k��}������☋��t�D��;��a�O��B�i�Q�n/#4'�Z�T���dY��C`������-�եf�ꍉ�qZ��#	�݊�cX�L�v����(u"�S4ƛhC���x:��D#�I���cLu)�r�v�=?�t�$�(�����/����f7�����^� Z��O�<ONe��cXj=G��H`w��1 ?���+�r�D�/^�y�景q���K��lr'a�
��������bѱT,`����#-��<* �x9�y�J��S�����Ar��ZR�J���RI'Z�JV��G�|/�:���И~� Ȳ� A/	(N�sA�N Є��a���yzB�k���"��T?��맛����|���u{gVsÌ39T����K�E��b���7��	�&��d�謮.����<���Rv�C�u�X;;�F�4�/���mȯ�%F^��'��#��j�%��<Ҩ��a���u�<a���-=i������+��O����H���1�F�0dmP�>N��b��d!2�ݎ���z���/^�1�Y~�Ce�p8j�y�RO����� 9t?qL�t��)�_�����l�D�[�B�S
��cy5�(�Z�X����L�Y��������T@���{��\=�U�2'��7�#*(0ӑ���>���i�ݽ��i*2::��{�ǭ�ނ�.�7N�^�aaaw��|�_�S��F��2��
�b��>��R����{��v	�1U��0��l��LvDӿmo"A5+�A���)Oڻ����� ��z��C�I����Jz&\
|�z�X�"  ��IDAT^������4>�֩��Q����z��Ɇ��d�Ml�<�lsO>|'J�y;�U�D�����E�b�B�n!'_�Е��ӲZ����\dHQ����Ƭ?\�hjLv˞	D�R4؊Y�Y��z��� @￸�q�cקK�F��GR�r�Nv
Tg@�h��<t�.�G��MW�#�������zTg�q|�M��Z�W�d"F9��D�r���x~�5�m��:=A�"���p���:�.����C(��V�v�'�.�B�o�
;}!��y矇믿�pllE.�ggg���O��{��������<Ǻ�!VǇd�m[7�����yу���uj�q���u^��>������'��<e%�-l�Ͳ��}&!l���_�D�uRo0)��1���ԧm�%�\�W���x��^�+��
##�v�K>_��%��Ën��;�1|������ V��8:x5��4(-"��&�S�2V�R�T��M����������Io����Vk��v�ǳ��C{ZX�x�j&>�>����Ԥ���9�5�o҉���(l�냯��eR��A0���ɛvm��8#���I�Cz�����2�g����߰KK2/A�o0����Qt�$��g���;*��JY�|�a\ZZ��Q�*����.�+�ӌ�Oƀ�ޏ����˪�{��.��F*���:ax����3<ZV(����<&:S���k���1?N��z!	��"�d �w{1�,��hf+yt˙�x4�J�/ade�i��q'(0~ᨴ3`�&p�[(�ɼ�mo����6\}��fg�ż����A�ڵ睷CCC�s�1?7ob�K��q����J����W�/�2��&��`���������xwSi�D�e��s�ՐJg0
k;�+�˹馛w���+p����q����}�{���2�S&)�+~�K�@�y�"��X����1�wKG*m���c=���z��0�vO&r�1� d��0��ߊ�n��������Z�x���?;t��?��Kx�t��IA2��0�|��Z>��cX�x��#�yp\j|Y�DM>�҉1m���m�r:v�<$w@��}�\�a�b,/}j��[�g{[z�lzӼ���mI��<�7�L~�e�� ����z:��:����R���q�	�������vs��:�$�9�}���1�A��R������k�x-��u��M�X�_�ھc;���Z��p�EG.)�8]��kC$NZ�`�A���A"�!�,�ΡdjB�'��R�����m�%��þ�.�s���`�F
\s�Ux���`[F7���OU"젎����?3_��s� �$}����ֆ(�
�Ifm]�e�D�Id��CO8��B̨;uY��tA	�T=|�a�?���{����a#i~n-pN'\d����Lz2��z��_��2�����ȏt����}���^F�Ǻ|�
��"z<��=[�Nl!Bd��������w�hM_.�o�.��N�}�k=�7��`�ۮ����R�^�	�-p�$"����ka��.*mu��z�/���	�75�#�ǚa?ֿ�#�y[�O�vz��	dw5?�.�l��� �h�Ӑ�"�5�y���
��]]�!�g�۶m�E]H� ���F�E���h�zS��weih y��Bx�TH+oj�L�C�G	zO�&�N�MNNbמ]�@�c�>+�{!y먿(���`b|��K6�%����$��%�:����:�dd�o�`�"�t#^�g�L�#Z�Awfg��H�lе�=m���	�������y��ͣI��krrz��v=z2����j<Z��)��ˣ��[0�:�����Ջ�&b�L�!�"�uz
���f>c��C���\��lNk���5e��i�y�������V�NK��4n�u�WGM{ך�ٖUj�\͕�\p�]d�f� �Z^���
&v�}�c��qBY���/;��J���kU�2��^[�vzE�y���9�<]LW~����D�˧1�n\rU.�'��{���e����RO�2S)qW�Hƣ��B��a�U�s�I4�U�x��ZJ#H�y㥃�בLD�tӥ���Y�"�ӯ��p|@8��$N�e�݁J�x��-�.|�A�0��H����2D���m�{[����m�͙��x�~�eX&��L��Ay��*�|�i��FM�!���h�[��|�+^ay��^���>!N��������ɍ�t�>:/�e��k�ͽ8c8���9(,&�q��J�	��Y�>�Z!��]��*�M��~�k�oߎ�[���l��hJ�+�&���@y��/�������U��@� ����e	\V�� Q�j=�n�ڠ.�&_U��0T��^��E%�@���B�����v�9��actc4��=[���l���|�i-rb�e�5:���X����"�۲��qPesK,-#[���c�P�`�NGT5'�h�ё����C����K�*�J5d�7�c�e��b�f�5]���8Fe (w+_B�4�2}�P{��u:�E�k�@Y��V���|��_���2�?�;��o{ı�#�+C���71nI�ERt���2g@4~�C%��g�����m�ӻmvJO���B]��3
b8��SC͎�Iź:O�̍���8F�a�0����y��t��\?�Ɖ:���#�_�D�?�X&R��Ѳ�\�Pq�����]�M�6�,�|W�r���ƍh���1��e��&Ok�����6������<v�����dR�`�����34R\�2�F��C�X	������K�i�$v�܁�����H��z������2,��B��� )���џ�e��|%;�,����փ"d�5����b>�s�ظ5��6�	�ZzY���Mf�:}��
�t���㵗��Ѩ��<~{�m/�|�6i`v��w�t7��I�v�8q�������c8rt/�|�q�&����3���زq?�������ĩ*�D7���{n���7	L��_u!n�p+�Z�4�@�+��a�~�vN����Ng�D��e;��7bq���y����⺭:�d2�����Á���Հw�nۃm���S,W[��M���ۮ݂�s8|�jtׯ�Ճ[�#莁�6�Б70{�S��K�m�\���ȟ��V�
Xr/]?Q ��4͍M���t���:h틘��,�J��F�G���XÚ�ƌm�Z��4�'�H��v��@��K޽��F	;*nu*��e�N��Ѫ���рG����rkѪ����OH�̢	���p��v�1�����Q�Iw85�1J�[��"�i�ӎ�խcL�G7l��aq1�
���p��I4[M?q�)��O�J#���>����x��$���8�Clsw\v.�<����!m�&�ق��_(>T!W�c#���R��xIqm�� *�v�:���2EaYC/oҦ;'�{��-�mY6 kEJ��f]��?m�(�X-���	�V�r5|�u%��[�bc	��|��x�U�x�yc�ެ�����F��6�-�nƻ�܈o�v�`;&Jl� ���Mx'�֑[Kx��y���q|���7n�ذ�3g�]{>�z�Fܾ;����q�8���Q\���N!��Y|����׎�;oډ��<���e[;xϋ���+ưg`ױ�������`hs�Vo�l?vp��[�ck�a��＼��^��t������s���L�5m1���7ޏ�O�'뷀�Zc~B�bm�
�	�O� 1l��؝Ȏ*d��L��dZfK��út�|�tD3zk�9Wx�ʲ�&�CiVV�CX�1�sFsG��<�t�4�a�O��,�h���'����ׄ-�w��XL��tAU$��(!��P�2��3��Gp1��L'����A'��a�P ^:�g�{v�
}2�D��S�VC�#�wOC�O?/��b���O{�5DH��'Bz�Е�� �k�<]���4����i��S�U���i�!�녮���)^v�m�r�F>��"K;v����	Ē6qC�u�)��I˭��:W
�_D���G�0�������U����B��;���z|������s������l��`��������-n�&f6;tC8or�.�4�|.�c�mLW�8�T����Cܕ�a����0��a�`K��la�<�Z9�k����U׋��x���xfj#�Q�r�lh�!����mj\tZf{��;���=����\ �mm���Z*ӏ�Ӻ�4�#:h"��'ZK{==F��+�I�F��ޏb�oGB�~��ql�Ms�!��t�kA̋�����D)0�/����#��eE���Ǐk���l�!p�� ���H����9����ti��Oή�[�y�l���>���CF�/��B�\{�vLV ~ʂ�f�)�)apZ�O89�J����ρG�]%�� I���Q��=����;�� ��[�Ǻ�a=X���A��jP����ֿ��+�-���j�u��v6���=QO�/���o���˧�܏������%��k6K���Y�<w�b�q�X	�m/�Qu.���|�8&�ػ�l��g��8R���"� ?[�i62x͋v ωWϖ0��g� 6�n6'<���L��z��%:���LlN��J����t.�kvepٶ"W��h�}R�Ѷ�M48���-LL)�0X?�y�eQN>���V��+?;
zxxJ_<�"!�>:Z��ޏi:K���G�G�p���`��k+!Q�3��HD�VN�djd���4�����KEX6�/��}yi䏇���5$�~:1��AH�y���	�dWح'�#p��xcN��h�n�$igqW*5��s��Xuw�� �eUK�.5vl�;Q������d�SY�9
S],�-]��HO��$�ɫFD�=u�֩����zf$���O0e& ����Փ��e�
T��-���P���2^�k���u���G�@$HF�$�ae���~�0�꽛q�XY:�;.�8w�2��M� s�(�QhȂ;T�w����B9\4��%[��1��2��G��`mE�z~m�����j���K�_�mv��n���C��<Z�%|��X;p��Ql�C۾1O�&�/4�T՟P5P�$.4ؒ��"�������l`%o�z/�����N<Xk�G�QIW6p5��D����Qz��|��(eq��R�c��L�U��T��.?"EZ5w�@���h�hl�1��J�ѱ��-���ԙ�xZƏ:�`a�3l�5L`�3L�6��Yt:��҅ƎPa���n��@Q8�n��zթ�1M��t����YѪ ���I��t���܌�E����G.|��M�"�a8�$�q�%�EY�M�tҨ/%�A��ɬt�Q�~�/o��'��%�([r�c8ͦ��,�8�Zb�V4�Nǌ>�u�Q�)u�j4�x�#6��9�F�y�Ԝ�gff����ꎘ���P{=�p~yT?NZ�U��p�0�nW���:8���}�Y�����/$�<���W��O|�Jj�֭���+�6Z{R<�`�gU��<"��˜8���1fh�O�U0���G��߾���)X�eQ&��ڌ�u?|�V��UW��m����9�i�ۛC3�������3��|�N5��ϠI��o���=�!ꡲ���B�Ω�cSU��-l(��&0��`j��/�LK��q�D�mЫ�280��j�����r�)C�\#���܁E��kw�e�m2�iw˱���[�Uʞ{`�̘+`x.K��g��8q�y�U�~-\�d/�!--��p�TtM��F�ꥰz���pR�½�_�zd]��q^���9�ej��T�"]<嗀��Y�
Abh�E�)��Sz$�{�崣�ڨ�oz����3��P]�������H]�Ӄ��/.,bzf�j��밗:CѮ�NGȼ��Sr&#!�kOqb3�1zF��*�����㏡V�ᡇ�n۹d�����j��~��R���vc���������ֵL0�%
	��e��.�E#W¥;'����l��n7p��al
�*
�&��y�U��n��ܶ�}��f���a-����q��<2�6vr�r�yc��νO��pWҬbG��kvq��B��N.���
tj��:�X������\�O,���A<��F��zɥ��kTN���fkXi�AC�'ղ�/�9l(-��^{�x�N�'�H�q��C`���kH:�\XAj�m@�7�iT�Z=笁ͷ�WT:��^H����ī�Z �~L�jϪ��J��^�c�ˤ�P9C��b$�71�6�i���G= �Be	m]E;���g5����i���̲A:�����2��#��d��8XW.f$�R��W�7��&�G��C=d��l�����4]ڸ����,Ӂg���-�ܺе��;�|?:�!"�&Z�F���@(�q�
��tZ�\������m8;;�G}���p-�襢'N���>����`R��;���Y�q�g��4G�%F�2,E�жHݽ��?��Ł�c?D��2v:�Sķ_�W�*`�|��<>��[�@oc��F�Ǉ��{z_����2���n2�b/���9��3l_�6`�ds�|���#�x�8w&Cy�d�c����z�;�<���4[X��MC�h�0Z�:L7
����(4�����0^ȡB�s��^DX�32v�6d��[��b5�����o���ON����*�t�M7I�
hp�b\��Kgf4���^p���u*��Z>I�h}B��`�=�����O���ʜ��.h��)��'�I�y���5Ғ�(����m�]����-���_@{��Q�(�T)}�°<[���~>�`s�Ǵ�>(��V�*e<�0��nvQ��g�A���j�@cڱ&0yM�7SV=���O|S��V����&,G#G%�|��q�f?wB:�ڭg-���l��R�8�4騘t������Wn�P<P�h\�-�b�]��������<�x�:#F���VO>�~���6�_��kf/�a�C�fm���#�V6��^N�~	ȇ�V%����}8���Y�p����S�$��O<��t�!A��t��7��i��o=������������Q�'���穻&�ut���:0>T@)����+8x�*�>r�:�2��ޠ�:���|�eo�=vj	��Aɯ�aq�YN���㾃8�����n����2k24�)6�8f
�c�؈=�z��ſ��3���8��i,��I�~�����U�Z�1#T��|P?�Ge�Xq��sW��o�hX��P>�Y�m�=9��d�8�C�H�V��i�:���R��EO�tKM��X&!��PaGU��#}�����xzIVC�}S�~��w}R�+�C�[�#�n���� I�� ү]�h���ıup��A����x�IƙuB����͙�9v��C?�&�d��<�rυ��X��I�qS�R��AT����;��;�u��x��/߅��{ s�h��"������?��x�J�'kL6���8l�����Du��=�ZA�4�Apn����W�<ʸhC��݄�۷�	��1=X�s�c��.�6��aώ��G�����H�tj����.��[x����P��'f����<��j��s�XY��S�UL�Ӊѡ����x��<e+��BϞ\�<n�1���BE7�4���W�-,�Z�
5~t��e{&��ہmc���TP�T0�k`�x���1�WNb�`�t�E6�*�?X��|"u�U$� ��F|��}�	�\]���!هg���ק<%�c�[;��g��/���	�]=
O������F#2�6��Y��&���Z�'ʾ
C�;�n�1��F� 6Ɗ�>�Ou�R��"�ӥ��'��9c���O�7�7��O~29�Sl���x��q7����?��.,-/���������ʹv�����{�ch1Ԙ��3������w��<l;�H�tU��]|Á&f�U�%��p].�y�&lذCC�hqվ��dJ���K�A�B.�o�ږ�	0.#�OR��x�Ƒ�:��IL7�`�`檍�� ��&`Z �q�e/�Lq3w9֩T��6�b�<�J����gȮ�u��Sx���<T���$�B��jܩ4�G���۟|��}x��v۴�[ a�;��NV�S��1��b��2��w_��wo��|��WO���b�D�[?�?z��x�[Qϔ��{���Ǳ��D�~�{_�7\<�:;��>w ���'1��dc
��;�C�nG3_�'��/���8N�w_�?�m��ı)��_���>�m;q�^�m�:z�n���:�������A|߫v��F��!Þ�.l93���[��>�v̫\Gk����@=��Һ�X�j�	:�x�럧�e��K�}�ŕ�#��x�����N��O�3����V�<I�ڙ��`j`R�g�,�����(��l��Bء7�ӕJ���>��m00�}��-�Y��劒�����L�&e�  X�i=�_�aP��$^?=`g����mw#Z�~��g6i��DC=�����zY�)/G�-��N��͋ǰc�9��*Eә�P��2�|?h��q	e���e�to���G�,���q���`�;��'�X�c�� ���?/m)3�#�[�v�U�/��1<����'�o7�ko���rw��܍�J�� �!ļs���Y�j���<�/r�����}��X'f$���A���f���s�D:�6�@qX�M^E�ޤ~qH�%P&�~�2]���IkwX�?��=��G��B���*u_��T��N���|�+M�-/aae3�*7꘩6i�s��lģs�xf�A�T����2E�J(�����م�Yi��
Ve�>�X��:�V�������tܩ�*t�9|����a<�r���b�+�J��9zϣ��D���:ej4��y7���'���,N�t@1p���weu���ۨQ���7K8VͣR]�|��Y�lk��V�OBx=Ј�?w��4�|�3%�4&BP`S��J�Z���a I �����(�~-�x��Z���Q�������ŶZms��R�3ڥ�Ꟍ{yKOן*�>��ڱFV��1�6g(G���w|z�j��p�`Uȡ��y�`��(�ʋ��P����Kל��t���s���ꃮ�\�.8_-+��
:պ�0��<� ���{�أ�ڵ�f�i�H��ޜ��M��Ӏ���:����ȃ��q�����ES�q�?ME���s�:���a?VdÃ���W���T�RB\��m��R�:��&ez�N��,�q;�J�ҩ����G�Q�[��FO�g�\��=3�'��(5�l�|�Wm��e�}Ά)�<ο�Ř-m	;��K��э���d�W%Eg}ms'�N+(�5Q�,��[�"�� �����al^�q;�j��g=���,�b��N��G�~�Kh�ǰ���ʢ�i`���N�$J:��v��(Wt��N��9j�QW��)4����X[F��ĝ�j��+lC#����	lhMs��1?��� �	А��0�����ip�S��C������/cn` ��u�6�9�3_��:Z(u*l� kM|��gP�}��N}��a#
�E<��|�Ko�֚�ec���
�#C	�k�����B1~��1{c��el6�h�ts���_��$��#�j�1r&��0��Xlșe�Ӽc{T_Vr�5}��+T�(!�<�|խ��&C�U���z��K�F�'�t���!�gM$���hߠ�a�F��;�o�&u��R��I�&��Ea�&��Ƃ0ߕ��
F��k�d�	�Ώխ�L����y,f|(�e�,��!�n�7�d}���a��Ȍ�=>W&�m\�{k��db��d�~�������|�&���X*��_�}]��{���lg��:��F�|Z��'q>�C�ӡ���⺙#*3�׮3X�����<^k2H�'��1p����J��l���ȁ�,��"�o%w���	ӻt~$���|n�q�v3��`�k@{gG��
a� 9Ń�i��7�Xo�Nb(�7��L �y���=��Z��A�&�n�h�}m�>�*�����1Q&�\��l�31>�:��b
��ɨi�kx��rԳ�c�n�D��eL׎��ևj��_����}0�9�A������D=(�ן6 �:���(����3^2��&4�=_�j�t���X��B�<�HX�� ��v:p�i�8�W"!�����FfY�W�l�`�ҭ�8����W%8�S8�d�������B5�29�g~����ă����.�t�y�z�Hw^f�ϕ�+��/Z�![�cAe�Nc�I�i�X?�Nœ��xИ`�W��zI��ǉZc-�jr\��n9A���x�m,rL���f���^���CvP��1H�u����/�iϒ�i��T^�!�P�x�o�5��\����:u�vx�-��'�x<_迡J�$���T�P��Ÿӱ#�<��ݖ�p��$6Z�U�:�`�� ��d��i�:��x�����├�,ׇ�S��NAB�o ֧S ]�������ǤH�8ȡD�#puu*^!1`�ju6�VF��q4��z8��43Ξn�*�v�sp�Χ��η�i�%�N{D�UҊ��+G����8�P~/�^� cN�W��|l����'���[g��~�(�a�GFT ��P�K�I��c��Pr$�`upr��5����\�F+���TG�GGӷ��̬#M��iR^�$տZ{�g�<;RV�����A��5�|gN�1�N�����:XO�����L�PZ�D�<a��On��]F�Y���26�ι��2RR������I����l����2���@�ɔ��A��L�L,4�l4N��&`ܡj��d��]vie˧0�*��dd������{��Sɒ��[O�B����(F&qr|��X�ʵ��Ʊ�oˋ��p"����l�V�AjNj�+�i������je�F������v`bA�m�q�}t���/��|byUʢ?>T�dZ�T�,PE��_��8�R:&��y��-��I����5����`G7�8�w>�
��浪��2*)}޸�sHM7�`���(�z�f�&�S���W� ������̶�X�����|v�_�KKۥ<;U���A����pK�0Q��ںQI[Gŋ�+p�Ulru���Y��¢��X�d��%�+DJ6�yT'5u����yLa-P�|�a�����`9=E/Ԅ�b���q<#h��)	��2�cJ:�/ &[V,ڇ���Zui�[B���n��������Z�!ČP����8�� �5��UD%�� mҩp |	�DZ�&�t�Q���.��Й@�]�pl�-�D��gϷ�$�Bk{D9U�n�l�Q����7�U�W�Q�-`�Q�ecC��	�5[��\%`;ru��6������Pn�8^[��u�w�V�B���.Y��R�X��d؝nԑ\"�F���WC�����9,/L!�x#�%LЀ�s�q�fyBG�i��H�d�2����6w�e��[�z�<ZX�T\��=��I��ld*j(]�,��wGJ�+��R�C�6O=�f1��xg�YL��K؊el��9�NaWq�Ju\@O���R���`�+�O�%�h�c��F�N't鉁�Q0������I�uk���{�	�Ǿ|r]/�
+Q��Q6V���� �.�>�!1D(dX�r���1�8MnoxR����F�G��������<,������sM4�49��h�Z�����8���wGr���Bc��A
3��������I���ɳN�PG��@%`5�4���:�����cK2U�^3����,�
�&L��k��H��\̓��s�D�5����Fۍl8)�d�+ח�.D���$�0W�sB���Y��(U��* :Jgi4t����.�Mn+GDcg���TŖL�:�:M:&�\�߇��҅�!7V���P���P�� �"?
��x8�n]�d�����H�YޚO0����6���`�OΧ�D��v���J��yd�fp�e�ڭ0Ѫ`���!·�l#�*q�X�Xg	��ʍ)��vx 珍�Xv�5*4�}��@S�4Ҳ���elh0hX%�U��2ת�T_Ba�r�3��]��Ӽb�V�M2G��a�a'i�.3M���f蔴�.��.���#� �j�sZ�j��N�$��OC˲ݥd��p��B�N;�����%,͜��[7���ak)��l�H��!�u�����rm�����F�cOn�q6�,AW��1�b[�b؀�;�F��ד�J��m���d�[T���bI�
e��M��B*M�O���K��R�t�<a7=K}�9�t
T�����bUHْ�Ma�6�%�ͱ���͸�����lr��J��o���
��ߺ�%=�!h��(X^M�H��w-�N�:.0���v�����p�il"�ܪ6�,P�q<��Uk�A�����Sz�
��ZuhKM��Ӏӛ<�S�*�ns֤�����L^���f�º��Tg(����"h�ׄJ����v�ǆV'F�S�#}�׀Tu^י��OH���,�N4ĕ�&�?1O���a1��F�i�ؗun���
Tߙ����.x"*���bNPr���m��"�H���*0��,W�'�r��94�Oa3w�s���]�0�H��RE�8��:W���+�C�����FR;���z{���[}�v8a�)����@�r�2@��N��4��e�
w�Or(����^&��>�e�-(�w܁���C�;=�d�nG�󻾔���	lY>�����.�8��+�l���&u��n��N�l�A]���W��ְel#y�&�ԫu�pj�G�b�+L[������e�E
y3Z��;�l�^�~]Pv�<���>Q�	�X�����{4rE�语j�(;���ȅ$�4�_;��z��i��n�G�zV�U���<FT�z��d��.�N_�Y;*,P?ə(N����@�X�]�������gPc�y\87MOU1'Th�#�b��R�hۮ����ʡ`J�� g@US2:��2�W9�W%��-��J�/7�LSDeT��H��Y����nl6?��ܠO,]'RM�\���v��1�z��fL�&��A�'��$NFEU������68y�&�t��rZ}���O�1�?�B� `�1���B���<��N���kiM�w��.X����~�GM�����'��_c�	Z�h�uH��a�����|���j����2�|r��hm�k.6�B�z��[E8Vi9����W����ϱƒ�[�wI�j�+#��nL�.Cg:\�vtG$%�s\�ݭtFz���ˮE!;���E���GƬ�L��#|�+^�W���غu+��#شy~��5�X��a�X���I��/���/�k��:a7�\~�Mȝw	���݋
��?O�>[���B���r8�^P��j�kdj�]V*vڰЬ�ݯ|)�r'��t���MZ0z��ZE�qWB�Z��?����_}�A�_���5��wG$R��n�Q�)�#� >�"W���4~=�o��"��0ȼ��)l\��"��rj�
��|�x���Q����#����v�u�.Ax��i���)���؊q����d=��`;�(����)���R�:�S��[�P�s>񆃝]��=��I���T�x��%nI��(sG�s�GuzR��c�#�<
cM$�'���Z)*�n����v�\h��� )h�k٢4�W���7^tɀ�x�V�iK��-���tA�Ogu��I���'�M��s>��^�<���&�`+�t�����)��!����ی���Ao�����8�oQ�&��"��v�������LkA�d\��ma;�~t>=w��9k�8��[t���d��#hr�E�����v��p׳����7m�+/߃|��q۩��F|l+����s��M���n-��7�7?�Y[�Jﮣ^��3c����q̩�-�l.հ�;�1��C�ì5�}=�Bv�~��������v3�O���x��^��;���;��޽{�3��gP����h"r���ذq��s��_���ɓ'��o��ݗ�O�� V��4����hK$���q��J���Ş֯VVР��j����꛱˘�-�]�呞uڥ 9���@go�R��7������e�﫼�4bY���F�n=����[�O-�o�z�R-��&�4hhm�@�83m�b^x�xW9cl�!�q��"BV�҉�S�V��Y'zE��;A���Uznx��$���Џ�(�_R��ϵ��c���G7�!SyJRy�I��ǩ� *��P��ġk�-ϐa�ѱ�����i���0��XɐG�lςTQ6T���
q�0�%ַ���6o�nd�+��7X��in�ȇ��]�
��;�My�u�;�k�~'�Xǆ�7��E4���?�ñ֠�{��H�E׺�ޖ�Q�mS�@σ�B���G�7�?���{��X��#��Gh�1K�.r:D�2d %�d�qD�Y.�
)ө0��М��?��v�! �\Go"2�:�D�t�o>���V�Ğ��z�L��o���/b��n��š�)�鿷�T�zj���>�w�Ǉ������ �����O}��6Ŝ�U�2.��2�?�y��pN凉#8\���B��E�Nfu]v���+�@M�ݭ��]���p�C*p'4��Ng��p��E���\I��Q���6�P��J=gtf��C}��O=�wQb]I����E��4�Ƌ�O_���ۉ�ԍ��/�ǰP�q��..*�<�"�K�1ڶ1��QںQ��QڻQں1���U�t�w�gp�2M���O��3���<6H�̌��������g�,���
��0N>e�����������|��s�ȃOr5�e'�m;(�NW'�QĖ&��;4�v]�Ut�6��qk )��*Oaylu%u��-�{��u�Έ��6����)8�ڊIa�l%��p��Nƫ��1�(�b�Ť�����I�Kf�܉
�d3�Hܐo<t�`N��]B�� 4~��ct!I��f��A:x/~����l�	�P���b	x��H
Lj�al`�����ANx�B#����`�j]#A�74�sވ{�Nmq�5j�J׊o�hC�E�S�`k�sm��J�L�0��"�J�Sh�`�9��ó�	<;5��( e2����-�ѥ���I)c0�M]����,q��P�'�0s�$r4ƃ�,�咊�����v:�z�+�k�N1�����>bz0��5��'��a|�C8��s9J�9��V2xvf�Ʃ@2:r񹞒Ya�˰r�Mbǌ?�x���M�p�ӡ��M?�}ŧ��p�1�>���a������b�s̏-Ob<���C���ݢa-��3�$3&$�aY؏�P�b�����Ck��O�v˽���2�~���ڰ�EUNy��,�RuY��z&�o��y��SȘ%�n��p�x$r���i������W��<�R�{��{p��1�]`�Q���R��#��ؿ+j�I�d�|E�׹Q��ʄn�M�C���;�:�����Y�I�
E-��V�r�|�&"%�����0A�"ĖV�=��8��0p��YA�7��	(����4x[���>_D��
���ծu��B��,��|�����"k�����qv��0>�po����0�l�x��x��n��K�;���!�~,�V���*���+�W��𝸰�9�_�vU¶
�g�Yd�S����Q'~A_�4Gu����J�R��;n���K�B	-�V�\i7�#lF��,ݞ�b�k�>�t��n�SO=�����w~睷��z��TVD�n�Tw�-w;�mK�!���ۭ�;J�6�{ƪ�� ��J%K�w�'��k�Ŗf1�x[�cc������!L�c�q���ۏͧ1�}�xǎ~+u:�L�vI\A�.teL�I�y.��ZЄO@�5dX�T�λ*��m���;:���Ŵx(义��kN��f�eϭ��/�&A�mY�ɥ��q#ᵋ��Q��:��v��똪�Ҝ*ќo�=��,2��W��@��"3�R�@��a���ݧ���q�ñ+��͢$��O{�Y$��?�v1+��aq�rv�AM5��Xч����G%I�y� �p ���z|�t�l@TgG��-H��@�����rH�ӫ�9$�|d��v}\��j;�w�̣�y�E��א1��
��.4i�k�8AV�q�߮q�T�ڃ,�|�b�=���,9/ڋ|A�6D#vfH�)����7,��)�݊
2U;��T��|>oo@���k�?������<y+��,��b���*���������tY'-�u-Ftf�"DY�i�A2�t$�v�ǲ�Ql5P @����*Y9f25�Y�2���6w�ܙz.��1G'Y�X��;�M���EϾt�\�e1MyS��~�jɕo�i�n<�o��<܅Dt�8�hs��4�8�]6I�
��p�e�U�`eEngu�:CǡW��(�҂@���ոug�FoП��--$c��C\�j(���m�W�}m���.�"h��v^;G�m%����l�P�K;��|ݖ����r��O~�$��u����)��4*��i���x�U ���6������4j4끉J���'�_�������a}���җi���軺y���?=�~�ר�Gc�ǂ���?V�z�d�7ϱ�F-��4�-?!��%��<~MF�"us��,���kӻ���� ��)��N���<ыD+�,�j�.�k��A�8~9ߘ�9,�A�.���~�'�ۿ������G�Ǘ�tju�
�z�'�x�xd�&癝�1�ex$c���͉��L2פO&_)�^fJ�6*ݏ]!�ߡ�i�2�C�t�\���&��
mk�s�s��W�ثf�o��3Jf��\7(̮�%��"�]�-��0��5�ׂ��f��.���v�o�VH����_�v�a�����t�@��89:u�T����I꺢�t1C�v�c�`6C�����1�Ԥ!o
kC�+Q �#k�~�_�O�9ZV�~�g���'O���ߏj�K�\�~�>��}�y�v<s�9��RP��e�b%6�ֽ�ߌۮڇ�O>��j�yE��_`î*W��{9~��w���o��J�p�yX�����*V�LCT|/�8�{��q�{03;�ٺ������݈7]{	FGp����k�W^�[�]���ۋ[/ڍ�/<7^x���3�hRA�2e����}}�NB�O�FgYlز+yݪ]tj��^F�hQ���c�aEg��g.P�W�'�7/�����1��B	�e]VjMR1obtp��C�|����fɨY��ك�%�/��蠶�C2���!ja�	��¨Uǋ6.c{���]N6eU���$�c�ɰNo��6��.͒|�nN�x�@����Z�F�g4id�� =�l�Q^��d�F�X�T�n��C�yt饗��/��;w�ċ^t���/�۰� �n\��V������e��\Uʹ�8W%��Mtҡ}TE82`�bD�A:��|dD[t&�ے��5+(Vȥh�լ�?�x)@׫���Q�8��)�;��nNb.#��a�3MZ�!�Q?Jہ$Mgy���]?�>HǸ^��m7_�w�H;w�v<��~.htIDh����^�c?��+q3m��Rs���;ně�ً޳�ˤo㖽c��ۮ�u�o��O<�JF�Or�Cߍ}��㯻���"����2-?���)������@c�@$���h��q���<*ͪ0S�k�C�:> |����n�
W�ނWB�";l���oz+��%��vazi�;!UX��&~���C��	�����ڭ�88�mƻ^t�㏿?��/��a������!|����{_q=vL�S���yz�W]�������K�`���U/ڇ���*���W���^�w��J����6*���۸�$GM�0��+��������ࠥ\��P�M�}��5i��'�Z�	�n���l��:3���^�$�pz�jc�&P/����A�RZMD�x3U.Ic,}ZX�U��ɘ�ѪS��5 �2H%�����ג"��������c�T����vV��+�Fq����1���N���$�wjj
�7oƖ-[��s����y>�m�#4y��n5�1S��>{;sغr[������ز��-�<Z�jn��Q<�AA����]�V�y����'jv u/�i8�kP�BE�ld��$SC�:��i���w�c�P��3r�΄�6��������/��_��v�ǈ�m����V���K�����\�g�i/�z���=�j�����e���W��w��;^}��l�uڑ��)`���x�V�����:>L]ƻ0�����}���"&v�~C�HbR�V<:�p�S�l�60��m�]��H��ʽ�wl�%;F96Z��}��Q󻿊�i����ï���2��u|����ݿ}��q_^Ħ�,��k����VlgX��w���?)9Oϫ#[d���7Ӷ5�w	����
.51��;��d���y쟣���׃N�����K�����+]��'�^\d���mՕ�4����C)Z��̍uN�`��
�����vFPܤ��L
׃��~��by<3�+���_�(k�<1]�P|a'K$a{�F�ӯ4cr<[�RH��7�NP���d��S���4��`t�$���~��s�t�w����KT<�&k�ݣj��ΔH_�P����c�=���(,���t�]z�c��F_�yzz
��ك�_����?��� �z����ɖr�}�Kpqyۚ'��q�M7������]��:�g�7>�b���&�f��^m��t��JL�]M��4�D�8�D�]��E)����ǂ	��g�>�5�ЪoM��Kr�,z������=�>��S���[^r#J��{+��O=$���ċ/ٍy<x�0����γ�1�E~���]OU��e������/�-[ȣ�E-3�]`E�R�'ݦNi�v���`;K!{�f�6�t�BJ��!m=m]�ǎ��=�Ls�
�~�^l/�Ӫ�"q۵b��J_y�)�=5���k�Ļ_y�ܩ���A��W�?�[�������c������{�'����0�	�A�B�vI��%Eq�i 2\��$�����#���:�ǧ�=�sl����_�'>�{�؝_A��]סb;�W*,��Ry��ZR����uȌ�WAL?��W�u��61��*d�"��QG�l�:�����i�݊0��R���s
�H��x!��=e�,N�P�n��j�v���+�-j=D^�ש��o5du�_;���}:�w�������7��ַ��:Ս�O���}Y9��-V�֝�ez�R�E��/yiqW$�^p� F^t�ʋ�t��J
$g��p��ӛ,l���H�dX�k:�
k�lmb��-Ț4�1:��S��=�h�s=M����[�p��q:ɨW��p�u�`5:���}?*da]i�:s>&�?��|�ko���2�ǃ�����)\�"�X�[��(��G�P�vB�����:�¢���G��4�i��7��ޗ������-�5<ud�9h;���n�����	�����{��١qT�큦'+��?�_��*���k/�����6��%�ɣS򘜴95QNH7�f���͜X����ܲ/fʘ�c%7�edsT[J�:oNe����ā�׾u�����6`CD�O_���Q�>�Zu�9���:��t����k0v����@��v2�r��|"#?�#�:yLU�'��完�O �
�k*GT6S�*��:v�O�>S��ߖ8[�k�qr`S�a�6x���8�Us�Ig�2�A<��j�7�ؾ�_�[6oA���._�K�K��ηJ��/=���x67�å��B_=>OCɕ�]��v��<j�3��ꂷ_�5����N�Q�;M�'�x)�'�d�N�Iϱ�fYk�!=L�ӀwaГ	�j��[��� �E���]���	51Z��Ƌ��L����������+xfj_98�F�@�űf�i˞��k�6���'�}��cXf�z�<T��Z�t#�}b_	\��\��������J1���� �������?��'V8Wkx�k��`FOd�q�h	l݄l��;����v�6nׇG0O'�'wދ�͢nhTs1Ъb��Y��_l��>}�Cؽi3vO�A/,RCzi��ܜ��IvBMVt�J����Xu[��+")�	fn9u���>,�oć�v�;�V�k,S:��L�-Q������jʔ>\'U����i��H��h㠵��Z��#Y�	�_r�����fj��:M:'���� ׷�,1A!���}��h�H҅i�lR�G7�k���c(�D�?IrB�l�6��H�a�`��ל��!v]@���nW�4pT��s|�V����5ݥ�a�&�ԜN��co��r}��mu*_|)_2Ft�<�c��7�����a�˭A�&174I�3�c\�>z|�>�$*�*�����糟�,�9�~��R�N������#CO���8Y��|��8��ln'f�/Ľe�w��յ%8���U�0<��^��5�huݵ�h{�$u�':����K�]'_���������=�+Tsx_�$���t�����Y���23�������
�.k�r��IlP;�l���8�m��|�0V(_��O��G�Mᘆ���c�c��/ڇ�/ڌv>�e��ʐ-��$7��h�]�"������v��&H/�=����W��<�O���@�Zzn�ZdR����C�3�'7�]��^|�E�Z�`�<�/>��(�Vlc��j�<V*̞��;_�*��z�����g�oc�<�mہj����\$�)&Nj"w=6w��:X�3А^��\{#�W����-ؔA�*O���j�`��v�2<�_�2���w�?Hֈ���j�kM�7C+������Ѩ�QYFfn�2+�r4�+'J�|��c��*��1�7�Ƙ��nt_-u�P�@d�[!OSRS�ú�J�S��1��x$%��Y�ӁM�t��Ö��ǵf�<yjo�k��"�Hf`�0W��燶��y�9�]�vaiq	��&q��a�ɟ���+-�dעXG�P@��Ce0�łN�c=���y�iN�p8�6�躋e���h���z���t\H:���Q���4�4*n].�m�-��d�]������� bo�ȳ��b�:�P	�؁M�y��u\v��`��j=s��Q���8��\O�em��>�yX��q��߈��o9_���l1D��3������Hu�Nc�f�x��m������ƞ��Z����$dj���KOpgSkc�����r��ㆫI0�{�cG��Kl}��|��^Q!� �t�<�|�[��l�$Z	� �"�$�&���?J��hbiI��S�l�p�/ڱ	/�|n�d3nٷ/�h78��\<U�\���e��&�9�����o&�:|���]���&��3�慖�v"�Gmժ�c��zK򶰈��^�c7o7�-ĭ#�eq�n�5��w��Eנ/�ev��@_{��-7���qH' '�7h�h�毣׫�}����:u���z��i�G��N�鬀�I�L��W�vgv��h��	d�s�N��mo����=����moE����(W���(� ������S�_����`��۱4��E�D�9Ȝ�(R���a:V�-�ha;-��})�6J3D�Rc+�, 쇞,*��_#�p:{P�=��Pc�]\�7�l�-���.�q��M(vjx��<r'�ݮ�$�%�A�c��f����-���y+�.ٵ�y�ؠ����N�ľn�x�E�p�%����6�o�pg��qn��>Ǎ��)O�[�œ�jjg��?��@���S��K/ݽ��r#�M�`�ÿ���ج�[��t��UE��02�aVRЖ�^���t>M�}���۷�@��:ϑK��t�M*D���S3Q���j��F������!O���Κa�ek-���������o��m��w�?��7b�N��z'^T գ��n��8�򵭸�L3E���Y��#�ѡ��i��C@�|{�i�e���wHڼN�1�������/f
���v��	��޻ʝ��
��%�r�?��Ģ5-e0Ρ7N��Lr+>\F���L���eC�l��{��\\=� ��`�^��mkڝ�6�<��$fW8�5����N��v�|Bg���N�MN�2�ds>�s99֥�^m:=��iљ8�8�G����OO����ٟ�����k��k����]�8��Fӏ���|���[�MY*捿^ӥ.Uok'�S8>��)��4&�KS��\_l�(��T���ln��o��
w�Ъh�u+���T<e�eg���)#�j���u0�0�>���\�vӍ}�^�I"�T�Ef'xTS���GC#�A�/S'�d��������0��+/�N=�+6�3��]���r��r�c�d2�W�ߝ��
����Ã�᪠�w\{5^y��V�?֭G^d��a��ko�/����w�x����܎!���Q�y�ܰ���D�.(��Cڕ�-Y2�[h����%��;_�J���C��p�c��ʩ�U�����)Z�b�[�7�x&�^n-�=U���k�*�dV����ȶ��kx��,G�*j����H~J�����I���丛)&0����KG�^-�W��V�p|SS�:5���Y�XT��	謌�J�%z�Tţ�-~�!�_8g�	�v7/h�N��'�	#��j��L��f��{�v/���/��|��s���}��8p��-v�4��BĸF?a����S�8BC8D��F5���8Vr�!�G�v��C�3�V˱����3�itn�ơ��,!~�$��x�*�_[����*��tZ��F��v^{!ʮzS5H�'O�3>���߇�����{��=v��	�i�(E��3u���l{�KVچFU:ܦn��ᒅ���x ���ہG%ٝ\�2��Q�S�1����˱�w\(^B�Ǵ�P:��X,�C܋�.dy��9&��9�P�}L��^�l@mPui� �%G�T�Gﺗ㢃퓣x���"拃��O�F�,���A��ĸl�"�M�9��?���qx�c�Y���&���՘��T�D����
fN-c~v	�s�[\B-[�E���fsyT�:��+A:dD��z ���_�� >��SXb�2.�:�<���'q�CH[v]��
��|���Q9N������w��%��i/n��qt��m�\��]w	wE���s8�Ԥ��b�F���魷n�dre]##�1ѧff\��!HP5D�2�F]WZ.��{w~?�;�?������g��_ٟV�)3����W~�x<dX8�Z���R�&�>?-��������&xl<[H��W.��:W�uw@M�|����±�148��oz�ݐ�{�.T�L�L[��-'���ӓ����D�w��[_Bcxfr��T�f/^��ql�%86p���O����7��+���/�b]�^��]�+�=�7B��:sP࢑�k���}���x��[������]�}۷c��zu��&X-�"��c�ƍ��;p�-�`����/��N�[�c:��PX���Ÿ.[Ņ�ǰ{�0��j��K�q���P�H���e{C����$U��ŰNß��
Ԇ/��q��>D'�\�ņ��7�`�&<���������U���Ō]��촎<���u4}���3)�����ubzYDc�S�!UT�g�0��>���f�h��v����f�رi�Q�27�ڙi������zо��e:��2���܇y�׎��uC��k�%����y~�?}�������_���1/"���֯���:���ڼ6T�N�m�>�!ӌN��Ux�-
����;��-�
��Buw�?�*W+�;m��}7X�>�y|l�st �w��J�����m�������_����o���~�oq	���/�Z�w��ћ>v��oߥUo݉w_5�_���a_�^��ҍ
�"k��F�N+Kg�w9i�f��R�r�ӵ:��px�������2�����r���]�24���m��J���*:�p�IZM��i�j��2,�G|>:�g�5`��|��1��h��/ �1ĝ���v�H~^'����g@F�v&ԥ���kG��jg��h/q�����a������x�[ތ|��w��%.�R궾L&%���m��4�
Ǣ�A`���p���x��b)7���(��߁����oé�pӉ:6a���v�Ş�,��%B�t4���gWh��Vs�B� =����?���8��}8��8���a���e��@iК�|Ā���&wG_����������9����}��T���>&��)��8�_q�����8���h8��&��*\����7z��.0���/)��T�NaZ~t�f�N��5_�Li+\�.��X��X�t����2W�K\�/�JX$��(��A{����t6una]�3���"d?��
�ƀ��/!m���}8ZX��hc�G-�e�5�����c+e(��R<3��^��:�
�ߟ�.�yԯ����m����^�v(���Z&�`=�w�:�O� �?x̵Y���&-B����ZO�2xz��gV2������6>U+22.=��e�ἱ	K�jc�yt�z2T��$�d��ҷ�_��.teh�.���SF��aM2�M�Y�In��ݟ|�}t�j�v�~������m��w|^s��(g顗�/~磸�Ђ��C��*�,~��?Jg�®�a����������.� u�ȏ�w>r -{�'�!'%��V�iFl���]my:#W�k;��\;�lC�r6
w1�[������_��R���Ӄ�"x?��ӳ�<j�	d��`�$w�PS]���G��ك�?���p�c��ڥ�X���&�$?�e�Ѱ����=��bZ�c�A;5B"���˸س�e Y�©[��w�r��	7}p�.[|��b��u�'3��xl���0���6?��+����؏��^l�t����_i�u��!�Eo$q]ː�-�/��u��*�~��Ӊ����V��W��L�Aa7�2��3M��G�麳���ѩL[Vh�Б�i�er�b
�pVz��Bv��\i���_֯�z��G�lfd2��k��a�.;��J+�q�}&���N9�ƅ~�VF�1����ר��b�2��v�:j�P�C�_j�F���^�{q:K���Ǿ�G�W�Z'm|�E=�P/��o���]�ƨe�� ֢	3�{.����ơaK���a
�ad̹&e�Lv���cxp�8.��E����kԛ`;�W9<|r?����o��r���+KV*8V+�?u/�ѯ�W|���B���b���<�?�G�O�O!_.�=ȕ	W1vσ���+E���}�r[�������v^��>Q������ci}�D#'��ˁuah~���@��j�2���7��.��K���?�Z�j�٨���/}�v>333�Ϝ��ԾN3y��C���c��Jc�q/�E��\Mg��cJr@zFM�ҹ$��| ���Ș��Qp/�a~����D�FhDO�6wu�<��/��qLg�p�^���s~{��\���T�hs*���i�Z�89�׽�ux׻���_������u�*`�Y�����X%�c�M8^܊��/������a(��Av����s9�p
��ہ�Իv�M�&���'� �� ��x�q��ozË�%�ِ<j�>&[wޛB8Q�!)�
lA���R!$CNۧ���9�G�p�;��=�ſ�!}-p���ת8���e{v��:�W��C�0�sN�V�&E����?�q���}j�P7��C�?��_WFRWt<��Us�!R��b���7>�O>;�-[��N��4妘\���čY��p@ie�R���Ɇ�Q8��_�`c���;��1<PF�ۿgO�`���\����"��N8��.[�=��-[0H�ǗN��B�A*i	�j��^X�h��]�N��p״�r�M�tb�"�cu$vL���\;7�R�ʉN�1AzН}�_x=�����V��ɀ���;���a�	��gz]�Iq��לh����:a]�H*]�c�,�#�X'�}W[6M�g��r�殦UYF}a�va���������]�صc'����wC������[��y��ǃBƖ�^�7��#o�Ѩ��G
j�EQ��7l��K��eһ��[�~&��i�l��I�U¾��}�|��ϱF�`Ic�"a�z�չV����@a�iu�Ս�G]R�4ѮVP��`ii˺�P]�԰e���G�u��8����P*1>>���Q8�쿘H�O�ei�'1=��;>:�\�6�dsLw�6������^�nT��C[4�|S��:c�����u�^� �Ί���.����#��2Y��0��_է��N�j�U[��|�=��~3�Ϛ���@rQ�S��5�Hl�5bE(�IQCzw��M��u��G��/�=#�b�e�s�#*{���r�y���C����b[��������(j$,�vqQ/k����l�@]�WJTo��9ne�T��&`?$*a�-�C�[�<nݻ	��=�b����>��4[U|��y<rr���Y�DⲜ.L�#�L�bg�n_�?���:I ei<��ѪNi���m��J���Ak,�g>;T��ق�a=�7�t"ē,wp��yz��V�z6@���%M�8Ý�����%A��{��5(m�8�(`�I4�[�B��%��&6��ɵى�Q�*�8g����i�f���l�Y�t�h���a�&5?	A?�R�
�0�e"��9nj�=�4�5�o^a��a��o�Swp��cjj��t{ы���wߍ�� 0�O�ҫ��t���_�_i��z��岜_����T���,�4*V��2�&��=C���O�p>�T2W�3�s//q���*w�1������ &���u�K*�h�����殝~��Q�z�s�\B]2S�c�
<T�1g\|ݦ@�����S��[�FgHG�f�7�Z���w����ޠ,��ӂ�G�''���ӥ�g��;/]������f�g���@����gã�D�:�B��� N�r8���׏�c�s�uhvSG���bߨM&��(��C*ny$!h��;�"Dz�%ZJ�m���y�e����6��Ҟ�!�ȹ/�?��ۄ���6SEn�,���کG���E���m��B���5v�o4&�Z��@}ꗓ�QJ(3��]q�%\�������~l���#h��;�L�Ĩ�'p�]hN��V[:���0��6=L��:�
M��+�h�t�P���r�HH� ���Aʠs�hs�g*�B�+x䑩�Zʢ-4g������+�_�+]"&ǀF�����s��Lle�����Z&��ȓ&����H�G�d�\����B�ս�қܷ(���ƨ�L����<�62L�����J�C�i���GQ�R0��*=�,>!ΟM�t�Vo#��7�}�h�;�:WqڙT1@�:��}��w(4D'O����C�7��Tm�ZM�\�8Z�ɑ�'��n�NG��2y:7�A�Pĩ�_�#3:���熆A��� qK�!��z%7���0�/��$wiZ��b��NN#�oU*���/�Hz��i��@{Y�>�s.Z�if7��玁X�����G���iٟ�i���=���,~�hd���+�ь�R%����H�ar(q�Jor�VyG���r��׮\B~I��n��)6KD'���PmP�e�l1M;1�c�`8��,�z���(��t3KC[���tZO�]Yg� SY�d2y��#�pT��q\j*؜'��QEZ�}���3�h�,� ���|f�PY�6�������ǮйPgԿ�W�SXY�u�7Y��D�_�Q�%[���m��kBl���t��N%�����q�.��/�V��������_����զ�M
�A���P�k4��t���V=^��*S��B;���Sg�3ӵPR�hs����Ԡ���4�(z�H:�t.W1��m��2v
Ĩ\*�n�]�lG�N�:�����Wi�'�@��;��Bq;'"��Դ�������"IU�E�]��8��	�m�/�M=�jm@��6T�.L�d<%!�����!Ms:H��¯='���L$У:��a�5��f8YNeTƬ��Q�m���g��;}�m܀Lc����գ�T8�V�-.bc��=�%��/��C?H��,�^�;v��/��_�Ħ-�]p>��W�ErNה�.�ߏ��f،
��Oep��}r�k��S3���t��"��n�x�T������g�lц4�~#7�c�'�IdcBQ�-�c�kfX�Q�t�:%��k(Թ��4,��H�\�I�P�E�B�eeF��N��P+a�0�:����i� �=�ʰƔ�KW�����͐��G�͞޵���W9����?'��[�i.'ÔOwV
�;��!#+�R&���>9e;FQ,=F���j����1^��$����y��Jʰ��Xٯ�d�0%� �Qk�o6Sa�#�98��qЯӓ��Hg��B�����؛����R��]/��;ƹ�7����y����O>9��!m��b��j��:5���dV�^=unMP��
ݱ8h��j���DLC���Yy��L��3�k�Ďq�P�*�p�S4^F��?�� ����S�[�߈��F�2��\}ق�!��O��/��>ň��)�5ְ�IAG��JXm1�� ����ř������\C��h��6� v�~(���#^�z����W���fL�`��7�n%�5%>N�6�|�R07�ҧm�-���	�
��X*���\�KM�6�N��؜����D�1T�X���,``��(WW���!<�ԓx��'�?����� 6mۉ����O���5��>-�M�ߧ��Ͱ��6hg���V�D9��K\�kk���{m���a׍�(QJ/���eZ�4L�HSҹ-"�:�J(m���5���C�,���d��i�6�k�UWN�D��i%���ks�c�.L���B&����o�Ƹ�%`DJT�s�*	��Y1;��sIcLvFq�6��4���
�ٰ���&�+���xT?���Ưi݃���2� qH��E��wD��4@ע@���b��7��S�� r�\�'-=��.lL�����z�a|�=��(�^��;�F�^$��'N����0�+Z�m�ϐTo�2�1�Њ�$3�,�_K�7�E+���	g@ԡ�0~�-�]������iY�)97������ke��b��L� `���S���N��Ķ�	�.4�ec/��f.V����Ǐ���¨iN��jؾ��o�k�qt�΂�^��B��O�D����c+�!L7G������喌��	��>�J=5 �eBװ3 >j'��f�k��T̏ ��Q����г�2~�ϏM�@#0����WT;�N_1R;h,�8���ˏt>$�����cn
��2:�%4*T�|v��t��8�|��U~�n�ްaK+Kؾk7��.������3bVCR�®W���M�xF��kz�|��堔��g�:�g^2^-3�L14�L�*��cjqD%�ދ)`�R$���h\9����Jj�igA#��&�n,��Q�n����*�J$���稰��&7�m�&�Vt\�y��Y��y�,�	J �Ȟ#�8��c��k������;YS`lE����-�=�չ~��V8���|���پu�5���Ǽ>A��d]YHkmU�1-�WO���T-Q���/�-�i��?�:�j�N���w���h�ܑ��Lvڒvp�����?��=�ȕ�����Ay;�Ÿ����i$�g�P�{W��J2A�QF��b�%�;%h�x��t������K���jQ���SZϩ��˧E���؎P|l�^\~׍Up�E�x��}���G_�������Q,nB'�Smu6�\r�~�~#��8	��%�LM���o���S�p�,/Wq�:�G+��.�A�]�Q�H,�Z�)���Q̷�+D�-$d��RM�cL��R�88E�ZJJ7	X�Ӥ�=�I�PJ�N]�P&�d�l�*����t�tXI������4�	�>��^�T����VЪUQY^���|��7a�+1�6#){eG���a<�|��,j���۪яz&�G�>���� Zɭ�H��ʰ��b��S��ۦk)L45�G���E����d���V�&D��d66B��c�jd�9ά�>�V�ȭbE�ӧ㱝u���cF):�U��&�ա�ٺd�J�Q�D���0`{;e
W,�|,�:�Ax���ӂ'��Gq�:/m�݆�a�Ă�X]/ �|�rQcԁzA���\�5��In�V���.L�[��s\�)Z`���/o�M��3�L~ن�6��*�5V�c��G�I�����O9�m ��ۇju�m]��k2��y:Ƶ��(�l�S�s2_��(~>t*:���N����,�����ӑQle����r~�|Y9-�]����Ņz��a�ʸP�z=I7��B1�
+��Ӆ�R�خr���'M��|����8?��p��<� S2��N��J󰕵רt����峌ǅMG:m����r������������Ƴ]���Q����>�TF�<����a�0���$:C�ȌlFt܈��$��XΑ�}k3�ݧ�	v�^]iÎ?��ўTTXƵ��},�]]Dݡ%̑^��ǫ��[Z��">Ə�Toॉ-~�6�
L��`F�Y2�4��A|C�X�N5��Y4��Aw~��=�9��S�(EC�|� ��"���B]�Q����d�ሶ�T�v���g��4���I��m6��k�˭���I�@e�K�k��:F̚�ZX��L&��g��%}�F�!�%=j�Q���\�hd��(���޵����;n{16���\��2Z#h����Ww.O�]G?�]����F�0�-�ƃ$�-Y(�e-��`l�`ExC� /�l,����/`C��l~aK�
�Є�=m�Hӏ���}�y��ꙑ=�UY�<y2��y�G�{�ϴ�Qq`��m��;B��K��f��g軻:)ex�X4*g4~���`�!ڵ��G��S��� �)���Z���pMY,L&��d�����#�4r�=w�,�eir m*O�D���b���&��'f�|sr��Ŀ�E�������qt��h2,�V�t��=׈���Z)����k��_<�w(��v) ���R�����x2���En�/�.��H]}<�q�-!�\ű{G�d�u3�<���u�D��	<��9d�*�V�� �����? mU���F[=t��m_��+��s�=��������
O	�m�?�L��s�{B�������X��k��F���+3����Xi�;ދ����n�� ��Wa�96�(�z8(�įr�W=0�����c-�㶡� ��O�(\R��>E3�d����B�LK8���Ȼ<!X}��{۲a��2�qNbpH1 l3.Z����8�B�(���\�ˋ���瞳D�?�0��x�����;��	���j-_��^6���v]���Wz}�z%�(�y��9n��v|��~�#���_v�V).�[��
��@��Dc�A�TNNeX3,��)#d �!(^�U�+0z7�4�i7�N3v1�3�t<��m2� b����L��D��VY�z��Ю��@;����	ޮw�H���@�`����i �"BNX w��"�u�Gq����Y�r�����V�&�e��@#�a� I�q?s-��x1�\n?��)�,l�}j?�%\D	�::u(}ج��|��ˈf�:���R�)�Q�`n}^������Yѿ��۾�5m���mO�[{��J��٥vZ�8'��y�� �ʛ���9� ���6B����A��n���:�͡��r+t<�Y(�ʐ�ޤw� D���GB��&ُ
3<[q�W��$��Ă��1�`g���6B�	>6o*?��T�a����}D�~�8:k̈Vh���+4�@�/T�.;���3�j�����s:��Δ�� iyA��|��|�=�������н�oG9��?.rsv@g� �;t�����k�/Fr��֏�E@�3�^��ȵ��^\���F31���t#��I,N[pt�Y�u�ЇIЄ�M��Þ��U�;��H@�{3Yp����ݼ��\�����wZ/8�tS�D��u��oWϡ}�*o�Gec�~r:i5�%ء�8��.���K�w�}1�aDv�#��:hn{�#,�m�e���޴����s�iIG��>J���Z���	ȕ��X�����	��U;��m?Q&(>H}CP�VgCD^�U�����?�^/G4����ﾚa眽`Y���I���mmP���c�]El����_6��u�M�7����r�EJ�6�7��2��l���W"c�E�ЛY�ka�#J�����v�D�C�S&{�8B�@i_k�2м�R� f�Δ�����A�nڮ:�V�̃l'�Xkm=n��!=Ӆ*�p��ny���;�׮X�m�;�([��jڶ��²�ſ2� ufX�z,��Xf�����q��ى�S4&.5:�v'�a�D�|��!�r��v��`p%�I,C�|��P�,~z�;$-6"�E��Bf�,�0�.�11!�L
jPk��sȘ�I��ÊGZ?�ĳ�0&���"e3/|��G����n�kрf�������ERqc��
)�|ʔ.�
ɬP���'��#	d�hp^?d��Z����\k��q�(>��pu
jG,��X��Q�*�h���G���%��D��6D[h�vdr�H���!�"z��y�KF�R�>h�1�~�iT�����������`W�硽����^J���\J��Ct]ӞB�����e*^��\ϸ�h�|c��l�:��]/+��z��D�����8/x#�m5�!,���R�+��UŲ\Kw�N����v|�\�����n9q�h����cf �����Cw���P���)�6ZA�%����5� �('Z׉����i*N4yr"r<a�i��\�2Ѐ�$�"ٙ�x���v��S"q�bB΁�D�ZqbmqAE �t�inKc�P1�ʌ�G�BNx��n���r��.�aKV�@�d^�Ac�t�\�ʁ�HG��`�tJ77I�]�,�4q^��hn/�5 _�.o�]W�5���WN+rCƺ�T��b�i0���?���8"yi��P���*��nq���Py�� ���B��z�C�i�H[h|�&�����)TB�t�C�I:����;��e�J�T�н���ȳ��'/b[4ap��:�>���>���d�e첑�A-����G��iO٩��8*�8�}�xȊ6�2E����������y�3�m� �t��dz\�]�ȆE��>�n �_�Pu���߬k}�i���^[��B?�l꼂ˏz��^|��r���=w���|���%3I<�|7ޥxş��ӭ����޾�ɇu$t���`d���j:Yuމ�3�}NTŠ������s�@�>�9��C�Nm)ʏ�)���H�Кxi���D2��Yic���	���a�I#3u�I;b�a,�t܌AR2r��R� �G���$�.p��Ǚ�Ko��nӬ8I���A��m��DΤ�O�!K2
ŗ�y�KN�/w�a�t}[�#=%T�DȻkx2��������Q!>!����ū�8m;
w�^��[=ϛ�ɴ� �c;�E�&~�x�S��6`�)+:h>�w}��/�+��?x��D<�I<�4Dh�Q��.���q{���������Ss
GPoЄ�_���ģE����z��_ǣlzL��d�r���#��Ǧ!Vٞ��q�r\�%Y���o���붹��?��~l��Y��-{�e[�mbG�ɛHY�ߘyQ��H@��AP��m�#W�M�hu4�U���5Ϲҝ��#/���k����pH�G�Pn����Y���!��	�9���ɉ����h<��ӫ�O����]�����-��j���1Lлc^I��>z�=�/���Wnyw[���Zsڶip&'Q'A�����.):8&è�p��1�|���3���披'E\����+��Ţ�;_C	�O.k��Ӹ#^�է�O��l�ܽ{�z 7�+��/���	�LB���/h�d���H%hq��$�'GEK
��;�mk#g��tf���u�5�UmnS�r�Ht2��̚L͜H�l�8�����]e0i�$!4	2���R�a�cr�|婅4�+?�g�&]^��U ���݁��DƝmܭ���(�o�a��'j��5�:��rӆt�o'��IT|�>��1���җ�������,S}�X:�'����N�K�H}��%�4�_x�|�Pv�taN����a<1>v�&-^�5Vّ��
i���a;��Ay�H=���m_���k#}�LFё-i�j\ѤٗerB_�	��[��z;��k<K��|Q�_��H��U��=�&E�����gT(ޢGA�Q?��.GXOv�r�-��Ô�c���?�/��AC��o�ၞ��CG2�;�<��Ⱥ����G9���܋������v���eDGű��s�:��66j���C1���Ջb	x�j;������?����m��*�h��| ��`IG(2g Iifnoo�h������7_�F{�ܸ��f��P\;A� �S����ME�� ��9R/L��5:1uU�q
 �:�?�Aw�!���䩂��s�LU˓����@;Rn�O>��h�b�X�I�g��kRؒ�Go|����v���v�ƃ���~Xu9�«����?��?���O�����>Ю�u�=��?j�_���s����k�O?�^:�\��]W��:�����߶nm�W�֢��V"J^�[ {v���ق%�/x? ��*��ʉ�Q���@�L��nHi�Ӌ�-h��Y%G�Zx��dG�`�p;��
AΥ���;��c%�Q\ R��.��ȗ�B'�H�쌚��	<�ѰӤw�߲%���R/�}���[Aԭ��X��x�{�eٶI�MG�e�*c��_�#Ζ��t&M�?)/(��xj�,��(Pz�ϖ؈�~�?�=zC� ����2Rݰ����>�	5� ��P�)y��JG<�Ρ?���^U��� �,L�:V!�e<}�!��an��$�r���)����PCݘ�qw�e1�-��v�8�Ά�1��.��ޱv�}�nh������l/s��� s@���}�Y�D�?�����=���O�o��O��?�l{ys�m�FmS��*�h�jPb�tn�ɉY�R�;��!�c~r�Q] �P�qJ��~�Y�y��d�s!"M94�ύg>:"v�"��5𙯵���i7ol��޸��練�R�q����}�ϵ�,>�b�]����q;|�*t-"+g��|���^=����;�ٖ6F�OM�?����_��h�������Ы���bt���y�@�R����_(mz@�h�{�1|�N��!zb2 �rCv�J�lC�V�0�F:���� �".MzHe��\N���|d66aO�7���PKl�� 30ǧ1YW	 �"W��$�����\O���J�0�;Wh�"��}0�����Fʓy�x��׋"z����/��r�!�1l� ۙ~ ���lJKv�F�j[��*^K!�"�v�w`��G$z}�6Q�A*Y���˻:��БL�d�F���	Z�	��o�O�<~K^@g��C�_��/8Ur�#��Ny�}��ș�	پ�G�!�o1�x=�Xs����v�5�hw_{U��ګ�{�s���j}�",��EpQ���Gp��и���I७������_�f����O{�ulljR��FJo�	���0h���o�1�o���~�ـm^��s7Q6� T"�]X��èr%;b��? ����l����t��������­kNj�y�7U�������#�cq�'�⳻ڮc����������������޻N�CG����j������{ڛ+�p�M�C��X�)�O1BL��j�!]�8�<~�&Y��JxEOu��>��>���tL��y}&����JG.�vq�w�.V�zN&�h��g������G~��j 70������~�mr��,�ݑ�NY��i�(�N?-�%���8'n��Ch&�v��s1��KT��[�܌S�\���3˪�A�v`>�d�]A�n Dr��>Tl��9�h��S����o;b�C�I��i�.��=�B�
F�a�z�v�����,����`N�H���*cK�%=<�+}
�ڰ�!�ə'�uy� ]�/�B�:�p!��e���C����7��ǿ>x�B�Q7�c�cm}�ݎ�O�=�]�>|�M�}G7ڱՑO��uБz�,�_}����J���(�-��<�w��~���^x����کN�ӯ��ξ�Ŕ���?e'���ΕQy=ahNv�������mN�A�p��s㫰�*�N%�tH�i�����R�P��{�}��v��W�闟i�Nn}��Ѓbi��#��+�T+���~�9�.W���Z|k�h��'�eGy�������Μ�]����U=wwd3G�����L�lldb�� >�B�`��p"�:�a���d�2��=��/U����P���w�kJ����Z!�:��0d(��	��PPt����Ɋ^�O�'���Y� ��<�x�ƅ�:�тV�����ŧ�OL�AؠA��#�pP�ya����'�������&�ڴ��t��<�*^|�q0�N��
k�PV0��1�+]�:~�/���=��!�f��!���7��թ�C�]����dz?�����j��uM�9�(���Ҏ>���([��c���Q;q�X;q�X�����G�CFmC���x-�r��}��9i����=��5�>9M�*Uy9"�Qyd�����sŇ�Eǈ(2KJ@e���3��Q�wAJw���oI�%�\G%u�pG���o�����o/��L�\�ϯ}Ⓝ�������q��(TN�����[��p��ȕ�.�����W���t��v��'��#+m���v��=�n��Ԭ|6�YM݈e�
8r�g *�C�����/���i���d!�R���B�WGn ��-0����Ű_�\�0���.	�ò"��� ��?�El &��'v.������m*��M>��"��=��R�v��#�K�6�^5�T�.(�i�r�<��C����?:{�.E�)�!��q&��p-���;��$�l8lB���>�#ٍ��%^8E��sf-��ɇIX�^�>q�G8���+C��$M!��Ah����Ɣ�`}���D8($�Dǂ�GA.�L����<Q~��͍�#me���p����6Y>'Q���V��J6u��T��]ΣJ�h�v/�[����>�Ik␱��{.���E�l�ȧ�F%B'>�[R�w��:XnfQ�_gR�EI[""5bB�����Q�ϡСx�C��C��h����W%���-�iUW��`�Q���󣄫_X�e'򱓆a�V�
Ү�7��P���9�]�lLܛ��2*�G#]"�ҳ(��AnV9�\�C.��=a$+V2�y�K�����r�r�8�-��u,����?w��B��)va�/�� t�q��,വ7�*�L����m~�O���    IEND�B`�PK   �]'Ut˩�  �"     jsons/user_defined.json�Ko�6�����Hp��ܶv��MI�=A���p$W�w��K9u܀vBK����iD}3��������7ݟ���Ɣq5]_��=A0�`���|X��<�?\e�õM[����UE�1wm�`WſYd��y��uiתTP�Wi�qjr� J������0�g�Ŧۚ� ��/�z�y��������w��u�\6U_<���~Y��U��hW�	cИB�]v8w�~۝#X��s�ۦ�gkCh.˛MW7wvۭh�z�S���(�XK�e"8�T��.��M�W�٫����r3�����l�ٻ�*[�>l���S.���O���=���W��ҁ�pp����s7� �Ů\��)���G.K��H.M9s���y
����î!�o��t���t��������t�[ e@�[!U@�[ft@��x:�,��G�dȔ�#�2dA�#�2d�b2m��k`T�����_�ǉoug;�'{�kצ�Ի�a��9�U"=p\^G7?^��r��@@���A-UѲ@���L�H30(+4�"er3a����)&������;�|��(I�T��K�1c���/h8������F����K�����|��r�ж�&��"\��WDT�Q��J#n�eJJ$�ІB����u�ð�����Q���!�&�vUDٶ*��6=�� ��#?�������{{�J�q��j���g�4E����%��KKD��\�\T��"�ޣ�28]^�����,Up�	P8�g������>��T�+�\{��V�׊Y�Y�Y�Y�Y���ڿ��Mvg���m�(�Ҵ4�mztU����*��ֹ$25��}�>]79���b��'��T��)��ҩ8����{�䷇�T�k��iK�A'L+L4S,�?8x���o�n��PK
   �]'U[?C8Gi  �0                  cirkitFile.jsonPK
   @'U��8nx;  �~  /             ti  images/21dc82dc-72ec-4a9d-931e-ac94256341be.jpgPK
   �K'Uu��@� �� /             9�  images/626defbd-9ffc-44de-b7fd-54699b7076eb.pngPK
   Y\"U8��Q�  > /             �F images/86525bf4-9941-42eb-811d-381dc5200b1d.jpgPK
   b^"U���3T  b�  /             d images/b0310726-02d1-40a2-b36d-0772497b5f9f.jpgPK
   9A'UD5�<� � /             �o images/bf05f532-b4f9-4ebd-a877-7859e21a15d5.pngPK
   �]'Ut˩�  �"               T jsons/user_defined.jsonPK      S  	   